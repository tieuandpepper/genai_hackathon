module lfsr(clk, rst, reinit, advance, out, initial_state, taps, out_state);
  wire _28_;
  wire _29_;
  wire _30_;
  wire _31_;
  wire _32_;
  wire _33_;
  wire _34_;
  wire _35_;
  wire _36_;
  wire _37_;
  wire _38_;
  wire _39_;
  wire _40_;
  wire _41_;
  wire _42_;
  wire _43_;
  wire _44_;
  wire _45_;
  wire _46_;
  wire _47_;
  wire _48_;
  wire _00_;
  wire _01_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  wire _08_;
  wire _09_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire _16_;
  wire _17_;
  wire _18_;
  wire _19_;
  wire _20_;
  wire _21_;
  wire _22_;
  wire _23_;
  wire _24_;
  wire _25_;
  wire _26_;
  wire _27_;
  input advance;
  wire advance;
  input clk;
  wire clk;
  input [4:0] initial_state;
  wire [4:0] initial_state;
  output out;
  reg out;
  output [4:0] out_state;
  wire [4:0] out_state;
  reg \out_state_reg[1] ;
  reg \out_state_reg[2] ;
  reg \out_state_reg[3] ;
  reg \out_state_reg[4] ;
  input reinit;
  wire reinit;
  input rst;
  wire rst;
  input [4:0] taps;
  wire [4:0] taps;
  assign _05_ = rst ? initial_state[0] : _27_;
  assign _28_ = _00_ ? 1'h0 : \out_state_reg[3] ;
  always_ff @(posedge clk)
    \out_state_reg[3]  <= _28_;
  assign _29_ = _00_ ? _03_ : \out_state_reg[2] ;
  always_ff @(posedge clk)
    \out_state_reg[2]  <= _29_;
  assign _30_ = _00_ ? _04_ : \out_state_reg[1] ;
  always_ff @(posedge clk)
    \out_state_reg[1]  <= _30_;
  assign _31_ = _00_ ? _05_ : out;
  always_ff @(posedge clk)
    out <= _31_;
  assign _06_ = rst | reinit;
  assign _00_ = advance | _06_;
  assign _32_ = initial_state[4] & _06_;
  assign _07_ = ~ _32_;
  assign _33_ = ~ _06_;
  assign _08_ = advance & _33_;
  assign _34_ = \out_state_reg[3]  & _08_;
  assign _09_ = ~ _34_;
  assign _35_ = _07_ & _09_;
  assign _01_ = ~ _35_;
  assign _36_ = initial_state[2] & _06_;
  assign _12_ = ~ _36_;
  assign _37_ = \out_state_reg[1]  & _08_;
  assign _13_ = ~ _37_;
  assign _38_ = _12_ & _13_;
  assign _39_ = _00_ ? _01_ : \out_state_reg[4] ;
  assign _03_ = ~ _38_;
  assign _40_ = initial_state[1] & _06_;
  assign _14_ = ~ _40_;
  assign _41_ = out & _08_;
  assign _15_ = ~ _41_;
  assign _42_ = _14_ & _15_;
  assign _04_ = ~ _42_;
  always_ff @(posedge clk)
    \out_state_reg[4]  <= _39_;
  assign _43_ = taps[0] & out;
  assign _16_ = ~ _43_;
  assign _17_ = taps[1] & \out_state_reg[1] ;
  assign _44_ = _16_ ^ _17_;
  assign _18_ = ~ _44_;
  assign _45_ = taps[2] & \out_state_reg[2] ;
  assign _19_ = ~ _45_;
  assign _20_ = taps[3] & \out_state_reg[3] ;
  assign _21_ = taps[4] & \out_state_reg[4] ;
  assign _46_ = _20_ ^ _21_;
  assign _22_ = ~ _46_;
  assign _47_ = _18_ ^ _22_;
  assign _23_ = ~ _47_;
  assign _24_ = reinit ? initial_state[0] : advance;
  assign _48_ = _19_ ^ _23_;
  assign _25_ = ~ _48_;
  assign _26_ = reinit | _25_;
  assign _27_ = _24_ & _26_;
  assign out_state = { \out_state_reg[4] , \out_state_reg[3] , \out_state_reg[2] , \out_state_reg[1] , out };
endmodule

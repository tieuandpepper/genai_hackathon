module counter(clk, rst, reinit, incr_valid, decr_valid, initial_value, incr, decr, value, value_next);
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  input clk;
  wire clk;
  input [1:0] decr;
  wire [1:0] decr;
  input decr_valid;
  wire decr_valid;
  input [1:0] incr;
  wire [1:0] incr;
  input incr_valid;
  wire incr_valid;
  input [3:0] initial_value;
  wire [3:0] initial_value;
  input reinit;
  wire reinit;
  input rst;
  wire rst;
  output [3:0] value;
  reg [3:0] value;
  output [3:0] value_next;
  wire [3:0] value_next;
  assign _064_ = _000_ ? _002_ : value[2];
  assign _065_ = value[3] ^ _030_;
  assign _037_ = ~ _065_;
  assign _066_ = _032_ ^ _037_;
  assign _038_ = ~ _066_;
  assign _039_ = reinit ? initial_value[3] : _038_;
  assign _067_ = ~ _039_;
  assign _040_ = _036_ | _067_;
  always_ff @(posedge clk)
    value[2] <= _064_;
  assign _041_ = _036_ & _039_;
  assign _042_ = _023_ | _025_;
  assign _068_ = _008_ & _011_;
  assign _043_ = ~ _068_;
  assign _044_ = _008_ | _011_;
  assign _069_ = ~ _018_;
  assign _045_ = _009_ | _069_;
  assign _070_ = _044_ & _045_;
  assign _046_ = ~ _070_;
  assign _071_ = _043_ & _046_;
  assign _047_ = ~ _071_;
  assign _072_ = ~ _047_;
  assign _048_ = _042_ & _072_;
  assign _073_ = _041_ & _048_;
  assign _049_ = ~ _073_;
  assign _050_ = _035_ | _049_;
  assign _074_ = _040_ & _050_;
  assign value_next[3] = ~ _074_;
  assign _075_ = _000_ ? _003_ : value[1];
  assign _051_ = _041_ & _047_;
  assign _076_ = _027_ & _051_;
  assign _052_ = ~ _076_;
  assign _053_ = _034_ & _052_;
  assign value_next[2] = _049_ ? _053_ : _035_;
  assign _077_ = _026_ & _041_;
  always_ff @(posedge clk)
    value[1] <= _075_;
  assign _054_ = ~ _077_;
  assign _055_ = _051_ ? _026_ : _054_;
  assign _078_ = _023_ ^ _055_;
  assign value_next[1] = ~ _078_;
  assign _079_ = _026_ ^ _041_;
  assign value_next[0] = ~ _079_;
  assign _080_ = rst | _007_;
  assign _056_ = ~ _080_;
  assign _081_ = value_next[3] & _056_;
  assign _057_ = ~ _081_;
  assign _082_ = rst & initial_value[3];
  assign _058_ = ~ _082_;
  assign _083_ = _057_ & _058_;
  assign _001_ = ~ _083_;
  assign _084_ = value_next[2] & _056_;
  assign _059_ = ~ _084_;
  assign _085_ = rst & initial_value[2];
  assign _060_ = ~ _085_;
  assign _086_ = _059_ & _060_;
  assign _002_ = ~ _086_;
  assign _087_ = _000_ ? _004_ : value[0];
  assign _088_ = value_next[1] & _056_;
  assign _061_ = ~ _088_;
  assign _089_ = rst & initial_value[1];
  assign _062_ = ~ _089_;
  assign _090_ = _061_ & _062_;
  assign _003_ = ~ _090_;
  always_ff @(posedge clk)
    value[0] <= _087_;
  assign _091_ = value_next[0] & _056_;
  assign _063_ = ~ _091_;
  assign _092_ = rst & initial_value[0];
  assign _005_ = ~ _092_;
  assign _093_ = _063_ & _005_;
  assign _004_ = ~ _093_;
  assign _094_ = incr_valid | decr_valid;
  assign _006_ = ~ _094_;
  assign _095_ = ~ reinit;
  assign _007_ = _006_ & _095_;
  assign _096_ = ~ _007_;
  assign _000_ = rst | _096_;
  assign _097_ = decr_valid & decr[1];
  assign _008_ = ~ _097_;
  assign _009_ = incr_valid & incr[0];
  assign _098_ = value[0] & _009_;
  assign _010_ = ~ _098_;
  assign _011_ = incr[1] & incr_valid;
  assign _099_ = value[1] & _011_;
  assign _012_ = ~ _099_;
  assign _100_ = value[1] ^ _011_;
  assign _013_ = ~ _100_;
  assign _014_ = _010_ | _013_;
  assign _015_ = _010_ ^ _013_;
  assign _101_ = _008_ & _015_;
  assign _016_ = ~ _101_;
  assign _017_ = _008_ ^ _015_;
  assign _018_ = decr_valid & decr[0];
  assign _102_ = value[0] ^ _009_;
  assign _019_ = ~ _102_;
  assign _103_ = _018_ & _019_;
  assign _104_ = _000_ ? _001_ : value[3];
  assign _020_ = ~ _103_;
  assign _105_ = _017_ & _020_;
  assign _021_ = ~ _105_;
  assign _023_ = reinit ? initial_value[1] : _017_;
  assign _106_ = _018_ ^ _019_;
  always_ff @(posedge clk)
    value[3] <= _104_;
  assign _024_ = ~ _106_;
  assign _025_ = reinit ? initial_value[0] : _024_;
  assign _026_ = ~ _025_;
  assign _107_ = _023_ & _025_;
  assign _027_ = ~ _107_;
  assign _028_ = _016_ & _021_;
  assign _108_ = _012_ & _014_;
  assign _029_ = ~ _108_;
  assign _030_ = value[2] & _029_;
  assign _031_ = value[2] ^ _029_;
  assign _109_ = ~ _031_;
  assign _032_ = _028_ & _109_;
  assign _033_ = _028_ ^ _031_;
  assign _034_ = reinit ? initial_value[2] : _033_;
  assign _035_ = ~ _034_;
  assign _110_ = ~ _027_;
  assign _036_ = _034_ | _110_;
endmodule

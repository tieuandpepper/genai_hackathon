module shift_left(out_valid, in, shift, fill, out);
  wire _192_;
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _025_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  input [11:0] fill;
  wire [11:0] fill;
  input [95:0] in;
  wire [95:0] in;
  output [95:0] out;
  wire [95:0] out;
  output out_valid;
  wire out_valid;
  input [2:0] shift;
  wire [2:0] shift;
  assign _003_ = shift[0] ? in[35] : in[47];
  assign out[89] = shift[2] ? _041_ : _038_;
  assign _042_ = shift[0] ? fill[8] : in[8];
  assign _043_ = shift[1] ? fill[8] : _042_;
  assign out[8] = shift[2] ? fill[8] : _043_;
  assign _044_ = shift[0] ? in[76] : in[88];
  assign _045_ = shift[0] ? in[52] : in[64];
  assign _046_ = shift[1] ? _045_ : _044_;
  assign _047_ = shift[0] ? in[28] : in[40];
  assign _048_ = shift[0] ? in[4] : in[16];
  assign _049_ = shift[1] ? _048_ : _047_;
  assign _004_ = shift[0] ? in[11] : in[23];
  assign out[88] = shift[2] ? _049_ : _046_;
  assign _050_ = shift[0] ? in[75] : in[87];
  assign _051_ = shift[0] ? in[51] : in[63];
  assign _052_ = shift[1] ? _051_ : _050_;
  assign _053_ = shift[0] ? in[27] : in[39];
  assign _054_ = shift[0] ? in[3] : in[15];
  assign _055_ = shift[1] ? _054_ : _053_;
  assign out[87] = shift[2] ? _055_ : _052_;
  assign _056_ = shift[0] ? in[74] : in[86];
  assign _057_ = shift[0] ? in[50] : in[62];
  assign _005_ = shift[1] ? _004_ : _003_;
  assign _058_ = shift[1] ? _057_ : _056_;
  assign _059_ = shift[0] ? in[26] : in[38];
  assign _060_ = shift[0] ? in[2] : in[14];
  assign _061_ = shift[1] ? _060_ : _059_;
  assign out[86] = shift[2] ? _061_ : _058_;
  assign _062_ = shift[0] ? in[73] : in[85];
  assign _063_ = shift[0] ? in[49] : in[61];
  assign _064_ = shift[1] ? _063_ : _062_;
  assign _065_ = shift[0] ? in[25] : in[37];
  assign _066_ = shift[0] ? in[1] : in[13];
  assign out[95] = shift[2] ? _005_ : _002_;
  assign _067_ = shift[1] ? _066_ : _065_;
  assign out[85] = shift[2] ? _067_ : _064_;
  assign _068_ = shift[0] ? in[72] : in[84];
  assign _069_ = shift[0] ? in[48] : in[60];
  assign _070_ = shift[1] ? _069_ : _068_;
  assign _071_ = shift[0] ? in[24] : in[36];
  assign _072_ = shift[0] ? in[0] : in[12];
  assign _073_ = shift[1] ? _072_ : _071_;
  assign out[84] = shift[2] ? _073_ : _070_;
  assign _074_ = shift[0] ? in[71] : in[83];
  assign _006_ = shift[0] ? in[82] : in[94];
  assign _075_ = shift[0] ? in[47] : in[59];
  assign _076_ = shift[1] ? _075_ : _074_;
  assign _077_ = shift[0] ? in[23] : in[35];
  assign _078_ = shift[0] ? fill[11] : in[11];
  assign _079_ = shift[1] ? _078_ : _077_;
  assign out[83] = shift[2] ? _079_ : _076_;
  assign _080_ = shift[0] ? in[70] : in[82];
  assign _081_ = shift[0] ? in[46] : in[58];
  assign _082_ = shift[1] ? _081_ : _080_;
  assign _083_ = shift[0] ? in[22] : in[34];
  assign _007_ = shift[0] ? in[58] : in[70];
  assign _084_ = shift[0] ? fill[10] : in[10];
  assign _085_ = shift[1] ? _084_ : _083_;
  assign out[82] = shift[2] ? _085_ : _082_;
  assign _086_ = shift[0] ? in[69] : in[81];
  assign _087_ = shift[0] ? in[45] : in[57];
  assign _088_ = shift[1] ? _087_ : _086_;
  assign _089_ = shift[0] ? in[21] : in[33];
  assign _090_ = shift[0] ? fill[9] : in[9];
  assign _091_ = shift[1] ? _090_ : _089_;
  assign out[81] = shift[2] ? _091_ : _088_;
  assign _008_ = shift[1] ? _007_ : _006_;
  assign _092_ = shift[0] ? in[68] : in[80];
  assign _093_ = shift[0] ? in[44] : in[56];
  assign _094_ = shift[1] ? _093_ : _092_;
  assign _095_ = shift[0] ? in[20] : in[32];
  assign _096_ = shift[1] ? _042_ : _095_;
  assign out[80] = shift[2] ? _096_ : _094_;
  assign _097_ = shift[0] ? in[67] : in[79];
  assign _098_ = shift[0] ? in[43] : in[55];
  assign _099_ = shift[1] ? _098_ : _097_;
  assign _100_ = shift[0] ? in[19] : in[31];
  assign _009_ = shift[0] ? in[34] : in[46];
  assign _101_ = shift[0] ? fill[7] : in[7];
  assign _102_ = shift[1] ? _101_ : _100_;
  assign out[79] = shift[2] ? _102_ : _099_;
  assign _103_ = shift[1] ? fill[7] : _101_;
  assign out[7] = shift[2] ? fill[7] : _103_;
  assign _104_ = shift[0] ? in[66] : in[78];
  assign _105_ = shift[0] ? in[42] : in[54];
  assign _106_ = shift[1] ? _105_ : _104_;
  assign _107_ = shift[0] ? in[18] : in[30];
  assign _108_ = shift[0] ? fill[6] : in[6];
  assign _010_ = shift[0] ? in[10] : in[22];
  assign _109_ = shift[1] ? _108_ : _107_;
  assign out[78] = shift[2] ? _109_ : _106_;
  assign _110_ = shift[0] ? in[65] : in[77];
  assign _111_ = shift[0] ? in[41] : in[53];
  assign _112_ = shift[1] ? _111_ : _110_;
  assign _113_ = shift[0] ? in[17] : in[29];
  assign _114_ = shift[0] ? fill[5] : in[5];
  assign _115_ = shift[1] ? _114_ : _113_;
  assign out[77] = shift[2] ? _115_ : _112_;
  assign _116_ = shift[0] ? in[64] : in[76];
  assign _011_ = shift[1] ? _010_ : _009_;
  assign _117_ = shift[0] ? in[40] : in[52];
  assign _118_ = shift[1] ? _117_ : _116_;
  assign _119_ = shift[0] ? in[16] : in[28];
  assign _120_ = shift[0] ? fill[4] : in[4];
  assign _121_ = shift[1] ? _120_ : _119_;
  assign out[76] = shift[2] ? _121_ : _118_;
  assign _122_ = shift[0] ? in[63] : in[75];
  assign _123_ = shift[0] ? in[39] : in[51];
  assign _124_ = shift[1] ? _123_ : _122_;
  assign _125_ = shift[0] ? in[15] : in[27];
  assign out[94] = shift[2] ? _011_ : _008_;
  assign _126_ = shift[0] ? fill[3] : in[3];
  assign _127_ = shift[1] ? _126_ : _125_;
  assign out[75] = shift[2] ? _127_ : _124_;
  assign _128_ = shift[0] ? in[62] : in[74];
  assign _129_ = shift[0] ? in[38] : in[50];
  assign _130_ = shift[1] ? _129_ : _128_;
  assign _131_ = shift[0] ? in[14] : in[26];
  assign _132_ = shift[0] ? fill[2] : in[2];
  assign _133_ = shift[1] ? _132_ : _131_;
  assign out[74] = shift[2] ? _133_ : _130_;
  assign _012_ = shift[0] ? in[81] : in[93];
  assign _134_ = shift[0] ? in[61] : in[73];
  assign _135_ = shift[0] ? in[37] : in[49];
  assign _136_ = shift[1] ? _135_ : _134_;
  assign _137_ = shift[0] ? in[13] : in[25];
  assign _138_ = shift[0] ? fill[1] : in[1];
  assign _139_ = shift[1] ? _138_ : _137_;
  assign out[73] = shift[2] ? _139_ : _136_;
  assign _140_ = shift[0] ? in[60] : in[72];
  assign _141_ = shift[0] ? in[36] : in[48];
  assign _142_ = shift[1] ? _141_ : _140_;
  assign _013_ = shift[0] ? in[57] : in[69];
  assign _143_ = shift[0] ? in[12] : in[24];
  assign _144_ = shift[0] ? fill[0] : in[0];
  assign _145_ = shift[1] ? _144_ : _143_;
  assign out[72] = shift[2] ? _145_ : _142_;
  assign _146_ = shift[1] ? _003_ : _001_;
  assign _147_ = shift[1] ? fill[11] : _004_;
  assign out[71] = shift[2] ? _147_ : _146_;
  assign _148_ = shift[1] ? _009_ : _007_;
  assign _149_ = shift[1] ? fill[10] : _010_;
  assign out[70] = shift[2] ? _149_ : _148_;
  assign _014_ = shift[1] ? _013_ : _012_;
  assign _150_ = shift[1] ? _015_ : _013_;
  assign _151_ = shift[1] ? fill[9] : _016_;
  assign out[69] = shift[2] ? _151_ : _150_;
  assign _152_ = shift[1] ? fill[6] : _108_;
  assign out[6] = shift[2] ? fill[6] : _152_;
  assign _153_ = shift[1] ? _021_ : _019_;
  assign _154_ = shift[1] ? fill[8] : _022_;
  assign out[68] = shift[2] ? _154_ : _153_;
  assign _155_ = shift[1] ? _027_ : _025_;
  assign _156_ = shift[1] ? fill[7] : _028_;
  assign _015_ = shift[0] ? in[33] : in[45];
  assign out[67] = shift[2] ? _156_ : _155_;
  assign _157_ = shift[1] ? _033_ : _031_;
  assign _158_ = shift[1] ? fill[6] : _034_;
  assign out[66] = shift[2] ? _158_ : _157_;
  assign _159_ = shift[1] ? _039_ : _037_;
  assign _160_ = shift[1] ? fill[5] : _040_;
  assign out[65] = shift[2] ? _160_ : _159_;
  assign _161_ = shift[1] ? _047_ : _045_;
  assign _162_ = shift[1] ? fill[4] : _048_;
  assign out[64] = shift[2] ? _162_ : _161_;
  assign _000_ = shift[0] ? in[83] : in[95];
  assign _016_ = shift[0] ? in[9] : in[21];
  assign _163_ = shift[1] ? _053_ : _051_;
  assign _164_ = shift[1] ? fill[3] : _054_;
  assign out[63] = shift[2] ? _164_ : _163_;
  assign _165_ = shift[1] ? _059_ : _057_;
  assign _166_ = shift[1] ? fill[2] : _060_;
  assign out[62] = shift[2] ? _166_ : _165_;
  assign _167_ = shift[1] ? _065_ : _063_;
  assign _168_ = shift[1] ? fill[1] : _066_;
  assign out[61] = shift[2] ? _168_ : _167_;
  assign _169_ = shift[1] ? _071_ : _069_;
  assign _017_ = shift[1] ? _016_ : _015_;
  assign _170_ = shift[1] ? fill[0] : _072_;
  assign out[60] = shift[2] ? _170_ : _169_;
  assign _171_ = shift[1] ? _077_ : _075_;
  assign _172_ = shift[1] ? fill[11] : _078_;
  assign out[59] = shift[2] ? _172_ : _171_;
  assign _173_ = shift[1] ? fill[5] : _114_;
  assign out[5] = shift[2] ? fill[5] : _173_;
  assign _174_ = shift[1] ? _083_ : _081_;
  assign _175_ = shift[1] ? fill[10] : _084_;
  assign out[58] = shift[2] ? _175_ : _174_;
  assign out[93] = shift[2] ? _017_ : _014_;
  assign _176_ = shift[1] ? _089_ : _087_;
  assign _177_ = shift[1] ? fill[9] : _090_;
  assign out[57] = shift[2] ? _177_ : _176_;
  assign _178_ = shift[1] ? _095_ : _093_;
  assign out[56] = shift[2] ? _043_ : _178_;
  assign _179_ = shift[1] ? _100_ : _098_;
  assign out[55] = shift[2] ? _103_ : _179_;
  assign _180_ = shift[1] ? _107_ : _105_;
  assign out[54] = shift[2] ? _152_ : _180_;
  assign _181_ = shift[1] ? _113_ : _111_;
  assign _018_ = shift[0] ? in[80] : in[92];
  assign out[53] = shift[2] ? _173_ : _181_;
  assign _182_ = shift[1] ? _119_ : _117_;
  assign _183_ = shift[1] ? fill[4] : _120_;
  assign out[52] = shift[2] ? _183_ : _182_;
  assign _184_ = shift[1] ? _125_ : _123_;
  assign _185_ = shift[1] ? fill[3] : _126_;
  assign out[51] = shift[2] ? _185_ : _184_;
  assign _186_ = shift[1] ? _131_ : _129_;
  assign _187_ = shift[1] ? fill[2] : _132_;
  assign out[50] = shift[2] ? _187_ : _186_;
  assign _019_ = shift[0] ? in[56] : in[68];
  assign _188_ = shift[1] ? _137_ : _135_;
  assign _189_ = shift[1] ? fill[1] : _138_;
  assign out[49] = shift[2] ? _189_ : _188_;
  assign out[4] = shift[2] ? fill[4] : _183_;
  assign _190_ = shift[1] ? _143_ : _141_;
  assign _191_ = shift[1] ? fill[0] : _144_;
  assign out[48] = shift[2] ? _191_ : _190_;
  assign out[47] = shift[2] ? fill[11] : _005_;
  assign out[46] = shift[2] ? fill[10] : _011_;
  assign out[45] = shift[2] ? fill[9] : _017_;
  assign _020_ = shift[1] ? _019_ : _018_;
  assign out[44] = shift[2] ? fill[8] : _023_;
  assign out[43] = shift[2] ? fill[7] : _029_;
  assign out[42] = shift[2] ? fill[6] : _035_;
  assign out[41] = shift[2] ? fill[5] : _041_;
  assign out[40] = shift[2] ? fill[4] : _049_;
  assign out[39] = shift[2] ? fill[3] : _055_;
  assign out[3] = shift[2] ? fill[3] : _185_;
  assign out[38] = shift[2] ? fill[2] : _061_;
  assign out[37] = shift[2] ? fill[1] : _067_;
  assign out[36] = shift[2] ? fill[0] : _073_;
  assign _021_ = shift[0] ? in[32] : in[44];
  assign out[35] = shift[2] ? fill[11] : _079_;
  assign out[34] = shift[2] ? fill[10] : _085_;
  assign out[33] = shift[2] ? fill[9] : _091_;
  assign out[32] = shift[2] ? fill[8] : _096_;
  assign out[31] = shift[2] ? fill[7] : _102_;
  assign out[30] = shift[2] ? fill[6] : _109_;
  assign out[29] = shift[2] ? fill[5] : _115_;
  assign out[2] = shift[2] ? fill[2] : _187_;
  assign out[28] = shift[2] ? fill[4] : _121_;
  assign out[27] = shift[2] ? fill[3] : _127_;
  assign _022_ = shift[0] ? in[8] : in[20];
  assign out[26] = shift[2] ? fill[2] : _133_;
  assign out[25] = shift[2] ? fill[1] : _139_;
  assign out[24] = shift[2] ? fill[0] : _145_;
  assign out[23] = shift[2] ? fill[11] : _147_;
  assign out[22] = shift[2] ? fill[10] : _149_;
  assign out[21] = shift[2] ? fill[9] : _151_;
  assign out[20] = shift[2] ? fill[8] : _154_;
  assign out[19] = shift[2] ? fill[7] : _156_;
  assign out[1] = shift[2] ? fill[1] : _189_;
  assign out[18] = shift[2] ? fill[6] : _158_;
  assign _023_ = shift[1] ? _022_ : _021_;
  assign out[17] = shift[2] ? fill[5] : _160_;
  assign out[16] = shift[2] ? fill[4] : _162_;
  assign out[15] = shift[2] ? fill[3] : _164_;
  assign out[14] = shift[2] ? fill[2] : _166_;
  assign out[13] = shift[2] ? fill[1] : _168_;
  assign out[12] = shift[2] ? fill[0] : _170_;
  assign out[11] = shift[2] ? fill[11] : _172_;
  assign out[10] = shift[2] ? fill[10] : _175_;
  assign out[9] = shift[2] ? fill[9] : _177_;
  assign out[0] = shift[2] ? fill[0] : _191_;
  assign out[92] = shift[2] ? _023_ : _020_;
  assign _192_ = shift[1] & shift[2];
  assign out_valid = ~ _192_;
  assign _001_ = shift[0] ? in[59] : in[71];
  assign _025_ = shift[0] ? in[55] : in[67];
  assign _027_ = shift[0] ? in[31] : in[43];
  assign _028_ = shift[0] ? in[7] : in[19];
  assign _029_ = shift[1] ? _028_ : _027_;
  assign out[91] = shift[2] ? _029_ : 1'h1;
  assign _030_ = shift[0] ? in[78] : in[90];
  assign _031_ = shift[0] ? in[54] : in[66];
  assign _032_ = shift[1] ? _031_ : _030_;
  assign _002_ = shift[1] ? _001_ : _000_;
  assign _033_ = shift[0] ? in[30] : in[42];
  assign _034_ = shift[0] ? in[6] : in[18];
  assign _035_ = shift[1] ? _034_ : _033_;
  assign out[90] = shift[2] ? _035_ : _032_;
  assign _036_ = shift[0] ? in[77] : in[89];
  assign _037_ = shift[0] ? in[53] : in[65];
  assign _038_ = shift[1] ? _037_ : _036_;
  assign _039_ = shift[0] ? in[29] : in[41];
  assign _040_ = shift[0] ? in[5] : in[17];
  assign _041_ = shift[1] ? _040_ : _039_;
endmodule

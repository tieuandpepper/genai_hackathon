module fifo_flops(clk, rst, push_ready, push_valid, pop_ready, pop_valid, full, full_next, empty, empty_next, push_data, pop_data, slots, slots_next, items, items_next);
  reg _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  reg _036_;
  reg _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_counter_items/value_loaden ;
  reg \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/gen_no_buffer.br_misc_unused_ram_rd_data_valid/unused ;
  wire \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/ram_rd_addr_update ;
  wire \br_fifo_ctrl_1r1w/bypass_ready ;
  wire \br_fifo_ctrl_1r1w/pop_beat ;
  wire \br_fifo_ctrl_1r1w/push_beat ;
  wire [7:0] \br_ram_flops/gen_read_data_pipe[0].br_ram_data_rd_pipe/gen_d[0].br_delay_valid_d/out_stages[0] ;
  reg [3:0] \br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] ;
  reg [3:0] \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] ;
  input clk;
  wire clk;
  output empty;
  wire empty;
  output empty_next;
  wire empty_next;
  output full;
  reg full;
  output full_next;
  wire full_next;
  output [3:0] items;
  wire [3:0] items;
  output [3:0] items_next;
  wire [3:0] items_next;
  output [7:0] pop_data;
  wire [7:0] pop_data;
  input pop_ready;
  wire pop_ready;
  output pop_valid;
  wire pop_valid;
  input [7:0] push_data;
  wire [7:0] push_data;
  output push_ready;
  wire push_ready;
  input push_valid;
  wire push_valid;
  input rst;
  wire rst;
  output [3:0] slots;
  wire [3:0] slots;
  output [3:0] slots_next;
  wire [3:0] slots_next;
  reg \slots_reg[1] ;
  reg [7:0] \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/mem  [12:0];
  always_ff @(posedge clk) begin
    if (_026_)
      \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/mem [\br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] ] <= push_data;
  end
  assign \br_ram_flops/gen_read_data_pipe[0].br_ram_data_rd_pipe/gen_d[0].br_delay_valid_d/out_stages[0]  = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/mem [\br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] ];
  assign items[3] = ~ _075_;
  assign _019_ = ~ _083_;
  assign _020_ = \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [0] & _026_;
  assign _021_ = \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [1] & _020_;
  assign _022_ = \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [2] & _021_;
  assign _023_ = \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [3] | _022_;
  assign _013_ = _019_ & _023_;
  assign _084_ = ~ _018_;
  assign _024_ = \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [2] & _084_;
  assign _014_ = _021_ ? _017_ : _024_;
  assign _015_ = \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [1] ^ _020_;
  assign _025_ = \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [0] ^ _026_;
  assign _016_ = _019_ & _025_;
  assign _085_ = \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_counter_items/value_loaden  ? full_next : full;
  assign _127_ = \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/ram_rd_addr_update  ? _000_ : \br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] [3];
  assign _086_ = rst ? 1'h0 : _085_;
  always_ff @(posedge clk)
    full <= _086_;
  assign _087_ = \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_counter_items/value_loaden  ? _028_ : items[1];
  assign _088_ = rst ? 1'h0 : _087_;
  reg \items_reg[1] ;
  always_ff @(posedge clk)
    \items_reg[1]  <= _088_;
  assign items[1] = \items_reg[1] ;
  assign _128_ = rst ? 1'h0 : _127_;
  assign _089_ = \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_counter_items/value_loaden  ? _029_ : items[0];
  assign _090_ = rst ? 1'h0 : _089_;
  reg \items_reg[0] ;
  always_ff @(posedge clk)
    \items_reg[0]  <= _090_;
  assign items[0] = \items_reg[0] ;
  assign _091_ = \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_counter_items/value_loaden  ? _030_ : _036_;
  assign _092_ = rst ? 1'h0 : _091_;
  always_ff @(posedge clk)
    _036_ <= _092_;
  always_ff @(posedge clk)
    \br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] [3] <= _128_;
  assign _093_ = \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_counter_items/value_loaden  ? _031_ : _037_;
  assign _094_ = rst ? 1'h0 : _093_;
  always_ff @(posedge clk)
    _037_ <= _094_;
  assign _095_ = \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_counter_items/value_loaden  ? _032_ : \slots_reg[1] ;
  assign _096_ = rst ? 1'h0 : _095_;
  always_ff @(posedge clk)
    \slots_reg[1]  <= _096_;
  assign _097_ = \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_counter_items/value_loaden  ? _033_ : \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/gen_no_buffer.br_misc_unused_ram_rd_data_valid/unused ;
  assign _098_ = rst ? 1'h0 : _097_;
  always_ff @(posedge clk)
    \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/gen_no_buffer.br_misc_unused_ram_rd_data_valid/unused  <= _098_;
  assign _099_ = \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_counter_items/value_loaden  ? _034_ : items[3];
  assign _100_ = rst ? 1'h0 : _099_;
  always_ff @(posedge clk)
    _075_ <= _100_;
  assign _101_ = \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_counter_items/value_loaden  ? _035_ : items[2];
  assign _102_ = rst ? 1'h0 : _101_;
  reg \items_reg[2] ;
  always_ff @(posedge clk)
    \items_reg[2]  <= _102_;
  assign items[2] = \items_reg[2] ;
  assign push_ready = ~ full;
  assign slots[0] = ~ items[0];
  assign slots[3] = ~ _036_;
  assign slots[2] = ~ _037_;
  assign empty = ~ \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/gen_no_buffer.br_misc_unused_ram_rd_data_valid/unused ;
  assign _129_ = \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/ram_rd_addr_update  ? _001_ : \br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] [2];
  assign \br_fifo_ctrl_1r1w/push_beat  = push_valid & push_ready;
  assign pop_valid = push_valid | \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/gen_no_buffer.br_misc_unused_ram_rd_data_valid/unused ;
  assign \br_fifo_ctrl_1r1w/pop_beat  = pop_ready & pop_valid;
  assign _064_ = slots[0] & \br_fifo_ctrl_1r1w/pop_beat ;
  assign _130_ = rst ? 1'h0 : _129_;
  assign _103_ = slots[0] ^ \br_fifo_ctrl_1r1w/pop_beat ;
  assign _065_ = ~ _103_;
  assign _066_ = \br_fifo_ctrl_1r1w/push_beat  & _065_;
  assign _067_ = \slots_reg[1]  & _064_;
  assign _104_ = \slots_reg[1]  ^ _064_;
  assign _068_ = ~ _104_;
  always_ff @(posedge clk)
    \br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] [2] <= _130_;
  assign _105_ = _066_ & _068_;
  assign _069_ = ~ _105_;
  assign _106_ = slots[2] & _067_;
  assign _070_ = ~ _106_;
  assign _107_ = _037_ ^ _067_;
  assign _071_ = ~ _107_;
  assign _072_ = _069_ | _071_;
  assign _073_ = _069_ & _071_;
  assign _108_ = _036_ & _070_;
  assign _074_ = ~ _108_;
  assign _109_ = slots[3] & _073_;
  assign _038_ = ~ _109_;
  assign _110_ = _066_ ^ _068_;
  assign _039_ = ~ _110_;
  assign _111_ = ~ _039_;
  assign _040_ = _038_ | _111_;
  assign _112_ = _073_ & _040_;
  assign _041_ = ~ _112_;
  assign _031_ = _072_ & _041_;
  assign slots_next[2] = ~ _031_;
  assign _042_ = _072_ & _074_;
  assign _113_ = _040_ & _042_;
  assign _030_ = ~ _113_;
  assign slots_next[3] = ~ _030_;
  assign _032_ = _038_ & _039_;
  assign _131_ = \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/ram_rd_addr_update  ? _002_ : \br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] [1];
  assign _043_ = items[0] & \br_fifo_ctrl_1r1w/push_beat ;
  assign _114_ = items[0] ^ \br_fifo_ctrl_1r1w/push_beat ;
  assign _044_ = ~ _114_;
  assign _045_ = \br_fifo_ctrl_1r1w/pop_beat  & _044_;
  assign _115_ = \br_fifo_ctrl_1r1w/pop_beat  ^ _044_;
  assign _029_ = ~ _115_;
  assign _132_ = rst ? 1'h0 : _131_;
  assign slots_next[0] = ~ _029_;
  assign _116_ = _032_ | slots_next[0];
  assign _046_ = ~ _116_;
  assign _047_ = _030_ & _046_;
  assign full_next = _031_ & _047_;
  always_ff @(posedge clk)
    \br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] [1] <= _132_;
  assign _048_ = items[1] & _043_;
  assign _117_ = items[1] ^ _043_;
  assign _049_ = ~ _117_;
  assign _118_ = _045_ & _049_;
  assign _050_ = ~ _118_;
  assign _051_ = _045_ | _049_;
  assign _119_ = _050_ & _051_;
  assign _052_ = ~ _119_;
  assign _053_ = items[2] & _048_;
  assign _120_ = items[2] ^ _048_;
  assign _054_ = ~ _120_;
  assign _121_ = ~ _054_;
  assign _055_ = _050_ & _121_;
  assign _056_ = items[3] | _053_;
  assign _122_ = items[3] & _055_;
  assign _057_ = ~ _122_;
  assign _028_ = _052_ & _057_;
  assign _058_ = _050_ | _121_;
  assign _059_ = _051_ | _057_;
  assign _123_ = _055_ & _059_;
  assign _060_ = ~ _123_;
  assign _124_ = _058_ & _060_;
  assign _035_ = ~ _124_;
  assign _061_ = _056_ & _059_;
  assign _133_ = \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/ram_rd_addr_update  ? _003_ : \br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] [0];
  assign _034_ = _058_ & _061_;
  assign _125_ = _028_ | _034_;
  assign _062_ = ~ _125_;
  assign _126_ = ~ _035_;
  assign _063_ = slots_next[0] & _126_;
  assign empty_next = _062_ & _063_;
  assign _134_ = rst ? 1'h0 : _133_;
  assign _033_ = ~ empty_next;
  assign \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_counter_items/value_loaden  = \br_fifo_ctrl_1r1w/push_beat  | \br_fifo_ctrl_1r1w/pop_beat ;
  assign pop_data[7] = \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/gen_no_buffer.br_misc_unused_ram_rd_data_valid/unused  ? \br_ram_flops/gen_read_data_pipe[0].br_ram_data_rd_pipe/gen_d[0].br_delay_valid_d/out_stages[0] [7] : push_data[7];
  assign pop_data[6] = \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/gen_no_buffer.br_misc_unused_ram_rd_data_valid/unused  ? \br_ram_flops/gen_read_data_pipe[0].br_ram_data_rd_pipe/gen_d[0].br_delay_valid_d/out_stages[0] [6] : push_data[6];
  always_ff @(posedge clk)
    \br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] [0] <= _134_;
  assign pop_data[5] = \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/gen_no_buffer.br_misc_unused_ram_rd_data_valid/unused  ? \br_ram_flops/gen_read_data_pipe[0].br_ram_data_rd_pipe/gen_d[0].br_delay_valid_d/out_stages[0] [5] : push_data[5];
  assign pop_data[4] = \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/gen_no_buffer.br_misc_unused_ram_rd_data_valid/unused  ? \br_ram_flops/gen_read_data_pipe[0].br_ram_data_rd_pipe/gen_d[0].br_delay_valid_d/out_stages[0] [4] : push_data[4];
  assign pop_data[3] = \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/gen_no_buffer.br_misc_unused_ram_rd_data_valid/unused  ? \br_ram_flops/gen_read_data_pipe[0].br_ram_data_rd_pipe/gen_d[0].br_delay_valid_d/out_stages[0] [3] : push_data[3];
  assign pop_data[2] = \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/gen_no_buffer.br_misc_unused_ram_rd_data_valid/unused  ? \br_ram_flops/gen_read_data_pipe[0].br_ram_data_rd_pipe/gen_d[0].br_delay_valid_d/out_stages[0] [2] : push_data[2];
  assign pop_data[1] = \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/gen_no_buffer.br_misc_unused_ram_rd_data_valid/unused  ? \br_ram_flops/gen_read_data_pipe[0].br_ram_data_rd_pipe/gen_d[0].br_delay_valid_d/out_stages[0] [1] : push_data[1];
  assign \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/ram_rd_addr_update  = \br_fifo_ctrl_1r1w/pop_beat  & \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/gen_no_buffer.br_misc_unused_ram_rd_data_valid/unused ;
  assign pop_data[0] = \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/gen_no_buffer.br_misc_unused_ram_rd_data_valid/unused  ? \br_ram_flops/gen_read_data_pipe[0].br_ram_data_rd_pipe/gen_d[0].br_delay_valid_d/out_stages[0] [0] : push_data[0];
  assign \br_fifo_ctrl_1r1w/bypass_ready  = pop_ready & empty;
  assign _004_ = \br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] [0] & \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/ram_rd_addr_update ;
  assign _005_ = \br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] [1] & _004_;
  assign _006_ = \br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] [2] & _005_;
  assign _007_ = \br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] [3] | _006_;
  assign _135_ = \br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] [2] ^ _005_;
  assign _008_ = ~ _135_;
  assign _002_ = \br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] [1] ^ _004_;
  assign _136_ = \br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] [0] ^ \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/ram_rd_addr_update ;
  assign _009_ = ~ _136_;
  assign _137_ = ~ _009_;
  assign _010_ = _002_ | _137_;
  assign _138_ = \br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] [3] & _010_;
  assign _011_ = ~ _138_;
  assign _012_ = _008_ | _011_;
  assign _000_ = _007_ & _012_;
  assign _139_ = ~ _008_;
  assign _001_ = _011_ & _139_;
  assign _003_ = _012_ & _137_;
  assign _140_ = _026_ ? _013_ : \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [3];
  assign _141_ = rst ? 1'h0 : _140_;
  always_ff @(posedge clk)
    \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [3] <= _141_;
  assign _076_ = _026_ ? _014_ : \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [2];
  assign _077_ = rst ? 1'h0 : _076_;
  always_ff @(posedge clk)
    \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [2] <= _077_;
  assign _078_ = _026_ ? _015_ : \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [1];
  assign _079_ = rst ? 1'h0 : _078_;
  always_ff @(posedge clk)
    \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [1] <= _079_;
  assign _080_ = _026_ ? _016_ : \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [0];
  assign _081_ = rst ? 1'h0 : _080_;
  always_ff @(posedge clk)
    \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [0] <= _081_;
  assign _017_ = ~ \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [2];
  assign _082_ = ~ \br_fifo_ctrl_1r1w/bypass_ready ;
  assign _026_ = \br_fifo_ctrl_1r1w/push_beat  & _082_;
  assign _018_ = \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [3] & _026_;
  assign _083_ = \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [2] & _018_;
  assign items_next = { _034_, _035_, _028_, _029_ };
  assign slots_next[1] = _032_;
  assign slots[1] = \slots_reg[1] ;
endmodule

module lfsr(clk, rst, reinit, advance, out, initial_state, taps, out_state);
  wire _28_;
  wire _29_;
  wire _30_;
  wire _31_;
  wire _32_;
  wire _33_;
  wire _34_;
  wire _35_;
  wire _36_;
  wire _37_;
  wire _38_;
  wire _39_;
  wire _40_;
  wire _41_;
  wire _42_;
  wire _43_;
  wire _44_;
  wire _45_;
  wire _46_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _09_;
  wire _11_;
  wire _13_;
  wire _15_;
  wire _16_;
  wire _17_;
  wire _18_;
  wire _19_;
  wire _20_;
  wire _21_;
  wire _22_;
  wire _23_;
  wire _24_;
  wire _25_;
  wire _26_;
  wire _27_;
  input advance;
  wire advance;
  input clk;
  wire clk;
  input [4:0] initial_state;
  wire [4:0] initial_state;
  output out;
  reg out;
  output [4:0] out_state;
  wire [4:0] out_state;
  reg \out_state_reg[1] ;
  reg \out_state_reg[2] ;
  reg \out_state_reg[3] ;
  reg \out_state_reg[4] ;
  input reinit;
  wire reinit;
  input rst;
  wire rst;
  input [4:0] taps;
  wire [4:0] taps;
  assign _05_ = rst ? initial_state[0] : _27_;
  assign _28_ = advance ? _02_ : \out_state_reg[3] ;
  always_ff @(posedge clk)
    \out_state_reg[3]  <= _28_;
  assign _29_ = advance ? _03_ : \out_state_reg[2] ;
  always_ff @(posedge clk)
    \out_state_reg[2]  <= _29_;
  assign _30_ = advance ? _04_ : \out_state_reg[1] ;
  always_ff @(posedge clk)
    \out_state_reg[1]  <= _30_;
  assign _31_ = advance ? _05_ : out;
  always_ff @(posedge clk)
    out <= _31_;
  assign _32_ = \out_state_reg[3]  & advance;
  assign _09_ = ~ _32_;
  assign _33_ = 1'h1 & _09_;
  assign _01_ = ~ _33_;
  assign _34_ = \out_state_reg[2]  & advance;
  assign _11_ = ~ _34_;
  assign _35_ = 1'h1 & _11_;
  assign _02_ = ~ _35_;
  assign _36_ = \out_state_reg[1]  & advance;
  assign _13_ = ~ _36_;
  assign _37_ = 1'h1 & _13_;
  assign _38_ = advance ? _01_ : \out_state_reg[4] ;
  assign _03_ = ~ _37_;
  assign _39_ = out & advance;
  assign _15_ = ~ _39_;
  assign _40_ = 1'h1 & _15_;
  assign _04_ = ~ _40_;
  always_ff @(posedge clk)
    \out_state_reg[4]  <= _38_;
  assign _41_ = taps[0] & out;
  assign _16_ = ~ _41_;
  assign _17_ = taps[1] & \out_state_reg[1] ;
  assign _42_ = _16_ ^ _17_;
  assign _18_ = ~ _42_;
  assign _43_ = taps[2] & \out_state_reg[2] ;
  assign _19_ = ~ _43_;
  assign _20_ = taps[3] & \out_state_reg[3] ;
  assign _21_ = taps[4] & \out_state_reg[4] ;
  assign _44_ = _20_ ^ _21_;
  assign _22_ = ~ _44_;
  assign _45_ = _18_ ^ _22_;
  assign _23_ = ~ _45_;
  assign _24_ = reinit ? initial_state[0] : advance;
  assign _46_ = _19_ ^ _23_;
  assign _25_ = ~ _46_;
  assign _26_ = reinit | _25_;
  assign _27_ = _24_ & _26_;
  assign out_state = { \out_state_reg[4] , \out_state_reg[3] , \out_state_reg[2] , \out_state_reg[1] , out };
endmodule

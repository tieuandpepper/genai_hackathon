module fifo_flops(clk, rst, push_ready, push_valid, pop_ready, pop_valid, full, full_next, empty, empty_next, push_data, pop_data, slots, slots_next, items, items_next);
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  reg _036_;
  reg _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  reg \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/gen_no_buffer.br_misc_unused_ram_rd_data_valid/unused ;
  wire \br_fifo_ctrl_1r1w/bypass_ready ;
  wire \br_fifo_ctrl_1r1w/push_beat ;
  wire [7:0] \br_ram_flops/gen_read_data_pipe[0].br_ram_data_rd_pipe/gen_d[0].br_delay_valid_d/out_stages[0] ;
  reg [3:0] \br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] ;
  reg [3:0] \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] ;
  input clk;
  wire clk;
  output empty;
  wire empty;
  output empty_next;
  wire empty_next;
  output full;
  reg full;
  output full_next;
  wire full_next;
  output [3:0] items;
  reg [3:0] items;
  output [3:0] items_next;
  wire [3:0] items_next;
  output [7:0] pop_data;
  wire [7:0] pop_data;
  input pop_ready;
  wire pop_ready;
  output pop_valid;
  wire pop_valid;
  input [7:0] push_data;
  wire [7:0] push_data;
  output push_ready;
  wire push_ready;
  input push_valid;
  wire push_valid;
  input rst;
  wire rst;
  output [3:0] slots;
  wire [3:0] slots;
  output [3:0] slots_next;
  wire [3:0] slots_next;
  reg \slots_reg[1] ;
  reg [7:0] \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/mem  [12:0];
  always_ff @(posedge clk) begin
    if (_026_)
      \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/mem [\br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] ] <= push_data;
  end
  assign \br_ram_flops/gen_read_data_pipe[0].br_ram_data_rd_pipe/gen_d[0].br_delay_valid_d/out_stages[0]  = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/mem [\br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] ];
  assign _019_ = ~ _082_;
  assign _020_ = \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [0] & _026_;
  assign _021_ = \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [1] & _020_;
  assign _022_ = \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [2] & _021_;
  assign _023_ = \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [3] | _022_;
  assign _013_ = _019_ & _023_;
  assign _083_ = ~ _018_;
  assign _024_ = \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [2] & _083_;
  assign _014_ = _021_ ? _017_ : _024_;
  assign _015_ = \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [1] ^ _020_;
  assign _025_ = \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [0] ^ _026_;
  assign _016_ = _019_ & _025_;
  assign _084_ = 1'h1 ? full_next : full;
  assign _124_ = \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/gen_no_buffer.br_misc_unused_ram_rd_data_valid/unused  ? _000_ : \br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] [3];
  assign _085_ = rst ? 1'h0 : _084_;
  always_ff @(posedge clk)
    full <= _085_;
  assign _086_ = 1'h1 ? _028_ : items[1];
  assign _087_ = rst ? 1'h0 : _086_;
  always_ff @(posedge clk)
    items[1] <= _087_;
  assign _125_ = rst ? 1'h0 : _124_;
  assign _088_ = 1'h1 ? _029_ : items[0];
  assign _089_ = rst ? 1'h0 : _088_;
  always_ff @(posedge clk)
    items[0] <= _089_;
  assign _090_ = 1'h1 ? _030_ : _036_;
  assign _091_ = rst ? 1'h0 : _090_;
  always_ff @(posedge clk)
    _036_ <= _091_;
  always_ff @(posedge clk)
    \br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] [3] <= _125_;
  assign _092_ = 1'h1 ? _031_ : _037_;
  assign _093_ = rst ? 1'h0 : _092_;
  always_ff @(posedge clk)
    _037_ <= _093_;
  assign _094_ = 1'h1 ? _032_ : \slots_reg[1] ;
  assign _095_ = rst ? 1'h0 : _094_;
  always_ff @(posedge clk)
    \slots_reg[1]  <= _095_;
  assign _096_ = 1'h1 ? _033_ : \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/gen_no_buffer.br_misc_unused_ram_rd_data_valid/unused ;
  assign _097_ = rst ? 1'h0 : _096_;
  always_ff @(posedge clk)
    \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/gen_no_buffer.br_misc_unused_ram_rd_data_valid/unused  <= _097_;
  assign _098_ = 1'h1 ? _034_ : items[3];
  assign _099_ = rst ? 1'h0 : _098_;
  always_ff @(posedge clk)
    items[3] <= _099_;
  assign _100_ = 1'h1 ? _035_ : items[2];
  assign _101_ = rst ? 1'h0 : _100_;
  always_ff @(posedge clk)
    items[2] <= _101_;
  assign push_ready = ~ full;
  assign _064_ = ~ items[0];
  assign slots[3] = ~ _036_;
  assign slots[2] = ~ _037_;
  assign empty = ~ \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/gen_no_buffer.br_misc_unused_ram_rd_data_valid/unused ;
  assign _126_ = \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/gen_no_buffer.br_misc_unused_ram_rd_data_valid/unused  ? _001_ : \br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] [2];
  assign \br_fifo_ctrl_1r1w/push_beat  = push_valid & push_ready;
  assign pop_valid = push_valid | \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/gen_no_buffer.br_misc_unused_ram_rd_data_valid/unused ;
  assign _127_ = rst ? 1'h0 : _126_;
  assign _066_ = \br_fifo_ctrl_1r1w/push_beat  & _064_;
  assign _067_ = \slots_reg[1]  & _064_;
  assign _102_ = \slots_reg[1]  ^ _064_;
  assign _068_ = ~ _102_;
  always_ff @(posedge clk)
    \br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] [2] <= _127_;
  assign _103_ = _066_ & _068_;
  assign _069_ = ~ _103_;
  assign _104_ = slots[2] & _067_;
  assign _070_ = ~ _104_;
  assign _105_ = _037_ ^ _067_;
  assign _071_ = ~ _105_;
  assign _072_ = _069_ | _071_;
  assign _073_ = _069_ & _071_;
  assign _106_ = _036_ & _070_;
  assign _074_ = ~ _106_;
  assign _107_ = slots[3] & _073_;
  assign _038_ = ~ _107_;
  assign _108_ = _066_ ^ _068_;
  assign _039_ = ~ _108_;
  assign _109_ = ~ _039_;
  assign _040_ = _038_ | _109_;
  assign _110_ = _073_ & _040_;
  assign _041_ = ~ _110_;
  assign _031_ = _072_ & _041_;
  assign slots_next[2] = ~ _031_;
  assign _042_ = _072_ & _074_;
  assign _111_ = _040_ & _042_;
  assign _030_ = ~ _111_;
  assign slots_next[3] = ~ _030_;
  assign _032_ = _038_ & _039_;
  assign _128_ = \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/gen_no_buffer.br_misc_unused_ram_rd_data_valid/unused  ? _002_ : \br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] [1];
  assign _043_ = items[0] & \br_fifo_ctrl_1r1w/push_beat ;
  assign _112_ = items[0] ^ \br_fifo_ctrl_1r1w/push_beat ;
  assign _029_ = ~ _112_;
  assign _129_ = rst ? 1'h0 : _128_;
  assign slots_next[0] = ~ _029_;
  assign _113_ = _032_ | slots_next[0];
  assign _046_ = ~ _113_;
  assign _047_ = _030_ & _046_;
  assign full_next = _031_ & _047_;
  always_ff @(posedge clk)
    \br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] [1] <= _129_;
  assign _048_ = items[1] & _043_;
  assign _114_ = items[1] ^ _043_;
  assign _049_ = ~ _114_;
  assign _115_ = _029_ & _049_;
  assign _050_ = ~ _115_;
  assign _051_ = _029_ | _049_;
  assign _116_ = _050_ & _051_;
  assign _052_ = ~ _116_;
  assign _053_ = items[2] & _048_;
  assign _117_ = items[2] ^ _048_;
  assign _054_ = ~ _117_;
  assign _118_ = ~ _054_;
  assign _055_ = _050_ & _118_;
  assign _056_ = items[3] | _053_;
  assign _119_ = items[3] & _055_;
  assign _057_ = ~ _119_;
  assign _028_ = _052_ & _057_;
  assign _058_ = _050_ | _118_;
  assign _059_ = _051_ | _057_;
  assign _120_ = _055_ & _059_;
  assign _060_ = ~ _120_;
  assign _121_ = _058_ & _060_;
  assign _035_ = ~ _121_;
  assign _061_ = _056_ & _059_;
  assign _130_ = \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/gen_no_buffer.br_misc_unused_ram_rd_data_valid/unused  ? _003_ : \br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] [0];
  assign _034_ = _058_ & _061_;
  assign _122_ = _028_ | _034_;
  assign _062_ = ~ _122_;
  assign _123_ = ~ _035_;
  assign _063_ = slots_next[0] & _123_;
  assign empty_next = _062_ & _063_;
  assign _131_ = rst ? 1'h0 : _130_;
  assign _033_ = ~ empty_next;
  assign pop_data[7] = \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/gen_no_buffer.br_misc_unused_ram_rd_data_valid/unused  ? \br_ram_flops/gen_read_data_pipe[0].br_ram_data_rd_pipe/gen_d[0].br_delay_valid_d/out_stages[0] [7] : push_data[7];
  assign pop_data[6] = \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/gen_no_buffer.br_misc_unused_ram_rd_data_valid/unused  ? \br_ram_flops/gen_read_data_pipe[0].br_ram_data_rd_pipe/gen_d[0].br_delay_valid_d/out_stages[0] [6] : push_data[6];
  always_ff @(posedge clk)
    \br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] [0] <= _131_;
  assign pop_data[5] = \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/gen_no_buffer.br_misc_unused_ram_rd_data_valid/unused  ? \br_ram_flops/gen_read_data_pipe[0].br_ram_data_rd_pipe/gen_d[0].br_delay_valid_d/out_stages[0] [5] : push_data[5];
  assign pop_data[4] = \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/gen_no_buffer.br_misc_unused_ram_rd_data_valid/unused  ? \br_ram_flops/gen_read_data_pipe[0].br_ram_data_rd_pipe/gen_d[0].br_delay_valid_d/out_stages[0] [4] : push_data[4];
  assign pop_data[3] = \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/gen_no_buffer.br_misc_unused_ram_rd_data_valid/unused  ? \br_ram_flops/gen_read_data_pipe[0].br_ram_data_rd_pipe/gen_d[0].br_delay_valid_d/out_stages[0] [3] : push_data[3];
  assign pop_data[2] = \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/gen_no_buffer.br_misc_unused_ram_rd_data_valid/unused  ? \br_ram_flops/gen_read_data_pipe[0].br_ram_data_rd_pipe/gen_d[0].br_delay_valid_d/out_stages[0] [2] : push_data[2];
  assign pop_data[1] = \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/gen_no_buffer.br_misc_unused_ram_rd_data_valid/unused  ? \br_ram_flops/gen_read_data_pipe[0].br_ram_data_rd_pipe/gen_d[0].br_delay_valid_d/out_stages[0] [1] : push_data[1];
  assign pop_data[0] = \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/gen_no_buffer.br_misc_unused_ram_rd_data_valid/unused  ? \br_ram_flops/gen_read_data_pipe[0].br_ram_data_rd_pipe/gen_d[0].br_delay_valid_d/out_stages[0] [0] : push_data[0];
  assign \br_fifo_ctrl_1r1w/bypass_ready  = pop_ready & empty;
  assign _004_ = \br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] [0] & \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/gen_no_buffer.br_misc_unused_ram_rd_data_valid/unused ;
  assign _005_ = \br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] [1] & _004_;
  assign _006_ = \br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] [2] & _005_;
  assign _007_ = \br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] [3] | _006_;
  assign _132_ = \br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] [2] ^ _005_;
  assign _008_ = ~ _132_;
  assign _002_ = \br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] [1] ^ _004_;
  assign _133_ = \br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] [0] ^ \br_fifo_ctrl_1r1w/br_fifo_pop_ctrl/br_fifo_pop_ctrl_core/gen_no_buffer.br_misc_unused_ram_rd_data_valid/unused ;
  assign _009_ = ~ _133_;
  assign _134_ = ~ _009_;
  assign _010_ = _002_ | _134_;
  assign _135_ = \br_ram_flops/gen_read_decoder[0].br_ram_addr_decoder_rd/gen_tiles_eq1.br_delay_valid_addr/out_stages[0] [3] & _010_;
  assign _011_ = ~ _135_;
  assign _012_ = _008_ | _011_;
  assign _000_ = _007_ & _012_;
  assign _136_ = ~ _008_;
  assign _001_ = _011_ & _136_;
  assign _003_ = _012_ & _134_;
  assign _137_ = _026_ ? _013_ : \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [3];
  assign _138_ = rst ? 1'h0 : _137_;
  always_ff @(posedge clk)
    \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [3] <= _138_;
  assign _075_ = _026_ ? _014_ : \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [2];
  assign _076_ = rst ? 1'h0 : _075_;
  always_ff @(posedge clk)
    \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [2] <= _076_;
  assign _077_ = _026_ ? _015_ : \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [1];
  assign _078_ = rst ? 1'h0 : _077_;
  always_ff @(posedge clk)
    \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [1] <= _078_;
  assign _079_ = _026_ ? _016_ : \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [0];
  assign _080_ = rst ? 1'h0 : _079_;
  always_ff @(posedge clk)
    \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [0] <= _080_;
  assign _017_ = ~ \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [2];
  assign _081_ = ~ \br_fifo_ctrl_1r1w/bypass_ready ;
  assign _026_ = \br_fifo_ctrl_1r1w/push_beat  & _081_;
  assign _018_ = \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [3] & _026_;
  assign _082_ = \br_ram_flops/gen_write_decoder[0].decoded_wr_addr[0] [2] & _018_;
  assign items_next = { _034_, _035_, _028_, _029_ };
  assign slots_next[1] = _032_;
  assign slots[1:0] = { \slots_reg[1] , _064_ };
endmodule

module tb;

    initial begin
        $display("TESTS PASSED");
        $finish;
    end

endmodule

module lfsr(clk, rst, reinit, advance, out, initial_state, taps, out_state);
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  wire _08_;
  wire _09_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire _16_;
  wire _17_;
  wire _18_;
  wire _19_;
  wire _20_;
  wire _21_;
  wire _22_;
  wire _23_;
  wire _24_;
  wire _25_;
  wire _26_;
  wire _27_;
  input advance;
  wire advance;
  input clk;
  wire clk;
  input [4:0] initial_state;
  wire [4:0] initial_state;
  output out;
  reg out;
  output [4:0] out_state;
  wire [4:0] out_state;
  reg \out_state_reg[1] ;
  reg \out_state_reg[2] ;
  reg \out_state_reg[3] ;
  reg \out_state_reg[4] ;
  input reinit;
  wire reinit;
  input rst;
  wire rst;
  input [4:0] taps;
  wire [4:0] taps;
  assign _028_ = ~ initial_state[4];
  assign _05_ = rst ? initial_state[0] : _27_;
  assign _029_ = _00_ ? _02_ : \out_state_reg[3] ;
  always_ff @(posedge clk)
    \out_state_reg[3]  <= _029_;
  assign _030_ = _00_ ? _03_ : \out_state_reg[2] ;
  always_ff @(posedge clk)
    \out_state_reg[2]  <= _030_;
  assign _031_ = _00_ ? _04_ : \out_state_reg[1] ;
  always_ff @(posedge clk)
    \out_state_reg[1]  <= _031_;
  assign _032_ = _00_ ? _05_ : out;
  always_ff @(posedge clk)
    out <= _032_;
  assign _06_ = rst | reinit;
  assign _00_ = advance | _06_;
  assign _033_ = _028_ & _06_;
  assign _07_ = ~ _033_;
  assign _034_ = ~ _06_;
  assign _08_ = advance & _034_;
  assign _035_ = \out_state_reg[3]  & _08_;
  assign _09_ = ~ _035_;
  assign _036_ = _07_ & _09_;
  assign _01_ = ~ _036_;
  assign _037_ = initial_state[3] & _06_;
  assign _10_ = ~ _037_;
  assign _038_ = \out_state_reg[2]  & _08_;
  assign _11_ = ~ _038_;
  assign _039_ = _10_ & _11_;
  assign _02_ = ~ _039_;
  assign _040_ = initial_state[2] & _06_;
  assign _12_ = ~ _040_;
  assign _041_ = \out_state_reg[1]  & _08_;
  assign _13_ = ~ _041_;
  assign _042_ = _12_ & _13_;
  assign _043_ = _00_ ? _01_ : \out_state_reg[4] ;
  assign _03_ = ~ _042_;
  assign _044_ = initial_state[1] & _06_;
  assign _14_ = ~ _044_;
  assign _045_ = out & _08_;
  assign _15_ = ~ _045_;
  assign _046_ = _14_ & _15_;
  assign _04_ = ~ _046_;
  always_ff @(posedge clk)
    \out_state_reg[4]  <= _043_;
  assign _047_ = taps[0] & out;
  assign _16_ = ~ _047_;
  assign _17_ = taps[1] & \out_state_reg[1] ;
  assign _048_ = _16_ ^ _17_;
  assign _18_ = ~ _048_;
  assign _049_ = taps[2] & \out_state_reg[2] ;
  assign _19_ = ~ _049_;
  assign _20_ = taps[3] & \out_state_reg[3] ;
  assign _21_ = taps[4] & \out_state_reg[4] ;
  assign _050_ = _20_ ^ _21_;
  assign _22_ = ~ _050_;
  assign _051_ = _18_ ^ _22_;
  assign _23_ = ~ _051_;
  assign _24_ = reinit ? initial_state[0] : advance;
  assign _052_ = _19_ ^ _23_;
  assign _25_ = ~ _052_;
  assign _26_ = reinit | _25_;
  assign _27_ = _24_ & _26_;
  assign out_state = { \out_state_reg[4] , \out_state_reg[3] , \out_state_reg[2] , \out_state_reg[1] , out };
endmodule

module enc_bin2onehot(clk, rst, in_valid, in, out);
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _00_;
  wire _01_;
  wire _02_;
  wire _05_;
  wire _07_;
  wire _08_;
  wire _09_;
  input clk;
  wire clk;
  input [3:0] in;
  wire [3:0] in;
  input in_valid;
  wire in_valid;
  output [14:0] out;
  wire [14:0] out;
  input rst;
  wire rst;
  assign _02_ = _01_ & _13_;
  assign out[1] = _00_ & _02_;
  assign out[0] = _00_ & 1'h0;
  assign _05_ = in[2] & in[3];
  assign out[14] = _05_ & 1'h0;
  assign out[13] = _02_ & _05_;
  assign out[12] = 1'h0 & _05_;
  assign _10_ = ~ in[2];
  assign _07_ = in[3] & _10_;
  assign _08_ = in[1] & _01_;
  assign out[11] = _07_ & _08_;
  assign out[10] = 1'h0 & _07_;
  assign _11_ = in[2] | in[3];
  assign out[9] = _02_ & _07_;
  assign out[8] = 1'h0 & _07_;
  assign _12_ = ~ in[3];
  assign _09_ = in[2] & _12_;
  assign out[7] = _08_ & _09_;
  assign _00_ = ~ _11_;
  assign out[6] = 1'h0 & _09_;
  assign out[5] = _02_ & _09_;
  assign out[4] = 1'h0 & _09_;
  assign out[3] = _00_ & _08_;
  assign out[2] = _00_ & 1'h0;
  assign _01_ = in_valid & in[0];
  assign _13_ = ~ in[1];
endmodule

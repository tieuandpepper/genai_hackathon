module cdc_fifo_flops_push_credit(push_clk, push_rst, pop_clk, pop_rst, push_sender_in_reset, push_receiver_in_reset, push_credit_stall, push_credit, push_valid, pop_ready, pop_valid, push_full, pop_empty, push_data, pop_data, push_slots, credit_initial_push, credit_withhold_push, credit_count_push, credit_available_push, pop_items
);
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  reg _0000_;
  reg _0001_;
  reg _0002_;
  reg _0003_;
  reg _0004_;
  reg _0005_;
  wire _0006_;
  reg _0007_;
  reg _0008_;
  reg _0009_;
  reg _0010_;
  reg _0011_;
  reg _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  reg _0048_;
  reg _0049_;
  reg _0050_;
  reg _0051_;
  reg _0052_;
  reg _0053_;
  reg _0054_;
  reg _0055_;
  reg _0056_;
  reg _0057_;
  reg _0058_;
  reg _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  reg _0069_;
  reg _0070_;
  reg _0071_;
  reg _0072_;
  reg _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  reg _0102_;
  wire _0103_;
  reg _0104_;
  wire _0105_;
  reg _0106_;
  wire _0107_;
  reg _0108_;
  reg _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  reg _0204_;
  reg _0205_;
  reg _0206_;
  reg _0207_;
  reg _0208_;
  reg _0209_;
  reg _0210_;
  reg _0211_;
  reg _0212_;
  reg _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  reg _0493_;
  reg _0494_;
  reg _0495_;
  reg _0496_;
  reg _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  reg _0528_;
  wire _0529_;
  reg _0530_;
  wire _0531_;
  reg _0532_;
  reg _0533_;
  wire _0534_;
  reg _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0541_;
  wire _0542_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0564_;
  wire _0565_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0572_;
  wire _0573_;
  wire _0575_;
  reg \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_bit_toggle_reset_active_push/src_bit_internal ;
  reg \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_gray_count_sync_push2pop/gen_cdc_sync[0].br_cdc_bit_toggle_inst/src_bit_internal ;
  reg \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_gray_count_sync_push2pop/gen_cdc_sync[1].br_cdc_bit_toggle_inst/src_bit_internal ;
  reg \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_gray_count_sync_push2pop/gen_cdc_sync[2].br_cdc_bit_toggle_inst/src_bit_internal ;
  reg \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_gray_count_sync_push2pop/gen_cdc_sync[3].br_cdc_bit_toggle_inst/src_bit_internal ;
  reg \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_gray_count_sync_push2pop/gen_cdc_sync[4].br_cdc_bit_toggle_inst/src_bit_internal ;
  reg \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_cdc_fifo_pop_flag_mgr/br_delay_nr_reset_active_pop/out_stages[1] ;
  wire [5:0] \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_cdc_fifo_pop_flag_mgr/push_count_adjusted ;
  reg [4:0] \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_cdc_fifo_pop_flag_mgr/push_count_saved ;
  wire \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_fifo_pop_ctrl_core/ram_rd_addr_update ;
  reg \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_gray_count_sync_pop2push/gen_cdc_sync[0].br_cdc_bit_toggle_inst/src_bit_internal ;
  reg \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_gray_count_sync_pop2push/gen_cdc_sync[1].br_cdc_bit_toggle_inst/src_bit_internal ;
  reg \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_gray_count_sync_pop2push/gen_cdc_sync[2].br_cdc_bit_toggle_inst/src_bit_internal ;
  reg \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_gray_count_sync_pop2push/gen_cdc_sync[3].br_cdc_bit_toggle_inst/src_bit_internal ;
  reg \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_gray_count_sync_pop2push/gen_cdc_sync[4].br_cdc_bit_toggle_inst/src_bit_internal ;
  reg [4:0] \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_saved ;
  wire [4:0] \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_visible ;
  wire [4:0] \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_credit_receiver/credit_incr ;
  wire \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/push_beat ;
  reg [7:0] \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][0] ;
  reg [7:0] \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][10] ;
  reg [7:0] \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][11] ;
  reg [7:0] \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][12] ;
  reg [7:0] \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][13] ;
  reg [7:0] \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][14] ;
  reg [7:0] \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][15] ;
  reg [7:0] \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][16] ;
  reg [7:0] \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][1] ;
  reg [7:0] \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][2] ;
  reg [7:0] \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][3] ;
  reg [7:0] \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][4] ;
  reg [7:0] \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][5] ;
  reg [7:0] \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][6] ;
  reg [7:0] \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][7] ;
  reg [7:0] \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][8] ;
  reg [7:0] \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][9] ;
  output [4:0] credit_available_push;
  wire [4:0] credit_available_push;
  output [4:0] credit_count_push;
  reg [4:0] credit_count_push;
  input [4:0] credit_initial_push;
  wire [4:0] credit_initial_push;
  input [4:0] credit_withhold_push;
  wire [4:0] credit_withhold_push;
  input pop_clk;
  wire pop_clk;
  output [7:0] pop_data;
  wire [7:0] pop_data;
  output pop_empty;
  wire pop_empty;
  output [4:0] pop_items;
  wire [4:0] pop_items;
  input pop_ready;
  wire pop_ready;
  input pop_rst;
  wire pop_rst;
  output pop_valid;
  wire pop_valid;
  input push_clk;
  wire push_clk;
  output push_credit;
  wire push_credit;
  input push_credit_stall;
  wire push_credit_stall;
  input [7:0] push_data;
  wire [7:0] push_data;
  output push_full;
  wire push_full;
  output push_receiver_in_reset;
  wire push_receiver_in_reset;
  input push_rst;
  wire push_rst;
  input push_sender_in_reset;
  wire push_sender_in_reset;
  output [4:0] push_slots;
  wire [4:0] push_slots;
  input push_valid;
  wire push_valid;
  assign _0554_ = ~ _0576_;
  assign _0577_ = _0035_ & _0036_;
  assign _0295_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][7] [6] | _0985_;
  assign _0296_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][3] [6] | _0208_;
  assign _0297_ = _0210_ & _0296_;
  assign _0578_ = _0295_ & _0297_;
  assign _0298_ = ~ _0578_;
  assign _0037_ = ~ _0577_;
  assign _0299_ = _0294_ & _0298_;
  assign _0300_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][4] [6] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][0] [6];
  assign _0579_ = ~ _0300_;
  assign _0301_ = _0210_ | _0579_;
  assign _0302_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][5] [6] | _0985_;
  assign _0303_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][1] [6] | _0208_;
  assign _0304_ = _0210_ & _0303_;
  assign _0580_ = _0302_ & _0304_;
  assign _0305_ = ~ _0580_;
  assign _0306_ = _0301_ & _0305_;
  assign _0581_ = _0035_ | _0036_;
  assign _0307_ = _0209_ ? _0299_ : _0306_;
  assign _0308_ = _0207_ | _0307_;
  assign _0582_ = _0290_ & _0308_;
  assign _0309_ = ~ _0582_;
  assign pop_data[6] = _0206_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][16] [6] : _0309_;
  assign _0038_ = ~ _0581_;
  assign _0310_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][13] [5] | _0985_;
  assign _0311_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][9] [5] | _0208_;
  assign _0312_ = _0210_ & _0311_;
  assign _0583_ = _0310_ & _0312_;
  assign _0313_ = ~ _0583_;
  assign _0314_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][12] [5] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][8] [5];
  assign _0315_ = _0314_ & _0988_;
  assign _0584_ = _0209_ | _0315_;
  assign _0316_ = ~ _0584_;
  assign _0585_ = _0313_ & _0316_;
  assign _0317_ = ~ _0585_;
  assign _0586_ = _0007_ | _0038_;
  assign _0318_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][14] [5] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][10] [5];
  assign _0587_ = ~ _0318_;
  assign _0319_ = _0210_ | _0587_;
  assign _0320_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][15] [5] | _0985_;
  assign _0321_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][11] [5] | _0208_;
  assign _0039_ = ~ _0586_;
  assign _0322_ = _0210_ & _0321_;
  assign _0588_ = _0320_ & _0322_;
  assign _0323_ = ~ _0588_;
  assign _0324_ = _0319_ & _0323_;
  assign _0589_ = _0209_ & _0324_;
  assign _0325_ = ~ _0589_;
  assign _0326_ = _0207_ & _0317_;
  assign _0590_ = _0325_ & _0326_;
  assign _0327_ = ~ _0590_;
  assign _0328_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][2] [5] | _0208_;
  assign _0591_ = ~ \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][6] [5];
  assign _0329_ = _0208_ & _0591_;
  assign \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_credit_receiver/credit_incr [4] = _0037_ & _0039_;
  assign _0592_ = _0210_ | _0329_;
  assign _0330_ = ~ _0592_;
  assign _0593_ = _0328_ & _0330_;
  assign _0331_ = ~ _0593_;
  assign _0332_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][7] [5] | _0985_;
  assign _0333_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][3] [5] | _0208_;
  assign _0334_ = _0210_ & _0333_;
  assign _0594_ = _0332_ & _0334_;
  assign _0335_ = ~ _0594_;
  assign _0336_ = _0331_ & _0335_;
  assign _0337_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][4] [5] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][0] [5];
  assign _0595_ = _0032_ | _0033_;
  assign _0596_ = ~ _0337_;
  assign _0338_ = _0210_ | _0596_;
  assign _0339_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][5] [5] | _0985_;
  assign _0340_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][1] [5] | _0208_;
  assign _0341_ = _0210_ & _0340_;
  assign _0040_ = ~ _0595_;
  assign _0597_ = _0339_ & _0341_;
  assign _0342_ = ~ _0597_;
  assign _0343_ = _0338_ & _0342_;
  assign _0344_ = _0209_ ? _0336_ : _0343_;
  assign _0345_ = _0207_ | _0344_;
  assign _0598_ = _0327_ & _0345_;
  assign _0346_ = ~ _0598_;
  assign pop_data[5] = _0206_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][16] [5] : _0346_;
  assign _0347_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][7] [4] | _0985_;
  assign _0348_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][3] [4] | _0208_;
  assign _0349_ = _0210_ & _0348_;
  assign _0599_ = _0007_ | _0040_;
  assign _0600_ = _0347_ & _0349_;
  assign _0350_ = ~ _0600_;
  assign _0351_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][6] [4] | _0985_;
  assign _0601_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][2] [4] | _0208_;
  assign _0352_ = ~ _0601_;
  assign _0041_ = ~ _0599_;
  assign _0602_ = _0210_ | _0352_;
  assign _0353_ = ~ _0602_;
  assign _0603_ = _0351_ & _0353_;
  assign _0354_ = ~ _0603_;
  assign _0604_ = _0350_ & _0354_;
  assign _0355_ = ~ _0604_;
  assign _0356_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][5] [4] | _0985_;
  assign _0357_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][1] [4] | _0208_;
  assign _0358_ = _0210_ & _0357_;
  assign _0605_ = _0356_ & _0358_;
  assign _0359_ = ~ _0605_;
  assign _0360_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][4] [4] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][0] [4];
  assign \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_credit_receiver/credit_incr [3] = _0034_ & _0041_;
  assign _0606_ = ~ _0360_;
  assign _0361_ = _0210_ | _0606_;
  assign _0607_ = _0359_ & _0361_;
  assign _0362_ = ~ _0607_;
  assign _0363_ = _0209_ ? _0355_ : _0362_;
  assign _0364_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][15] [4] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][11] [4];
  assign _0365_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][13] [4] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][9] [4];
  assign _0366_ = _0209_ ? _0364_ : _0365_;
  assign _0367_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][14] [4] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][10] [4];
  assign _0368_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][12] [4] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][8] [4];
  assign _0369_ = _0209_ ? _0367_ : _0368_;
  assign _0042_ = _0029_ & _0030_;
  assign _0370_ = _0210_ ? _0366_ : _0369_;
  assign _0371_ = _0207_ ? _0370_ : _0363_;
  assign pop_data[4] = _0206_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][16] [4] : _0371_;
  assign _0372_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][6] [3] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][2] [3];
  assign _0373_ = _0210_ | _0372_;
  always_ff @(posedge push_clk)
    _0001_ <= \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_gray_count_sync_pop2push/gen_cdc_sync[0].br_cdc_bit_toggle_inst/src_bit_internal ;
  assign _0374_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][7] [3] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][3] [3];
  assign _0608_ = ~ _0374_;
  assign _0375_ = _0210_ & _0608_;
  assign _0609_ = _0207_ | _0375_;
  assign _0376_ = ~ _0609_;
  assign _0610_ = _0373_ & _0376_;
  assign _0611_ = _0007_ | _0042_;
  assign _0377_ = ~ _0610_;
  assign _0378_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][11] [3] | _0208_;
  assign _0379_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][15] [3] | _0985_;
  assign _0380_ = _0210_ & _0379_;
  assign _0612_ = _0378_ & _0380_;
  assign _0013_ = ~ _0611_;
  assign _0381_ = ~ _0612_;
  assign _0382_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][14] [3] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][10] [3];
  assign _0613_ = ~ _0382_;
  assign _0383_ = _0210_ | _0613_;
  assign _0614_ = _0381_ & _0383_;
  assign _0384_ = ~ _0614_;
  assign _0615_ = _0207_ & _0384_;
  assign _0385_ = ~ _0615_;
  assign _0616_ = _0377_ & _0385_;
  assign _0386_ = ~ _0616_;
  assign _0387_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][13] [3] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][9] [3];
  assign _0388_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][5] [3] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][1] [3];
  assign \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_credit_receiver/credit_incr [2] = _0031_ & _0013_;
  assign _0389_ = _0207_ ? _0387_ : _0388_;
  assign _0390_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][12] [3] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][8] [3];
  assign _0391_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][4] [3] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][0] [3];
  assign _0392_ = _0207_ ? _0390_ : _0391_;
  assign _0393_ = _0210_ ? _0389_ : _0392_;
  assign _0394_ = _0209_ ? _0386_ : _0393_;
  assign pop_data[3] = _0206_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][16] [3] : _0394_;
  assign _0395_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][13] [2] | _0985_;
  assign _0396_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][9] [2] | _0208_;
  assign _0397_ = _0210_ & _0396_;
  assign _0014_ = _0024_ & _0027_;
  assign _0617_ = _0395_ & _0397_;
  assign _0398_ = ~ _0617_;
  assign _0399_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][12] [2] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][8] [2];
  assign _0400_ = _0399_ & _0988_;
  assign _0618_ = _0209_ | _0400_;
  assign _0401_ = ~ _0618_;
  assign _0619_ = _0398_ & _0401_;
  assign _0402_ = ~ _0619_;
  assign _0403_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][14] [2] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][10] [2];
  assign _0620_ = ~ _0403_;
  assign _0404_ = _0210_ | _0620_;
  assign _0621_ = _0007_ | _0014_;
  assign _0405_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][15] [2] | _0985_;
  assign _0406_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][11] [2] | _0208_;
  assign _0407_ = _0210_ & _0406_;
  assign _0622_ = _0405_ & _0407_;
  assign _0408_ = ~ _0622_;
  assign _0015_ = ~ _0621_;
  assign _0409_ = _0404_ & _0408_;
  assign _0623_ = _0209_ & _0409_;
  assign _0410_ = ~ _0623_;
  assign _0411_ = _0207_ & _0402_;
  assign _0624_ = _0410_ & _0411_;
  assign _0412_ = ~ _0624_;
  assign _0413_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][2] [2] | _0208_;
  assign _0625_ = ~ \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][6] [2];
  assign _0414_ = _0208_ & _0625_;
  assign _0626_ = _0210_ | _0414_;
  assign _0415_ = ~ _0626_;
  assign _0627_ = _0413_ & _0415_;
  assign _0416_ = ~ _0627_;
  assign \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_credit_receiver/credit_incr [1] = _0028_ & _0015_;
  assign _0417_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][7] [2] | _0985_;
  assign _0418_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][3] [2] | _0208_;
  assign _0419_ = _0210_ & _0418_;
  assign _0628_ = _0417_ & _0419_;
  assign _0420_ = ~ _0628_;
  assign _0421_ = _0416_ & _0420_;
  assign _0422_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][4] [2] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][0] [2];
  assign _0629_ = ~ _0422_;
  assign _0423_ = _0210_ | _0629_;
  assign _0424_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][5] [2] | _0985_;
  assign _0630_ = _0043_ ^ _0025_;
  assign _0425_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][1] [2] | _0208_;
  assign _0426_ = _0210_ & _0425_;
  assign _0631_ = _0424_ & _0426_;
  assign _0427_ = ~ _0631_;
  assign _0428_ = _0423_ & _0427_;
  assign _0016_ = ~ _0630_;
  assign _0429_ = _0209_ ? _0421_ : _0428_;
  assign _0430_ = _0207_ | _0429_;
  assign _0632_ = _0412_ & _0430_;
  assign _0431_ = ~ _0632_;
  assign pop_data[2] = _0206_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][16] [2] : _0431_;
  assign _0432_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][6] [1] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][2] [1];
  assign _0433_ = _0210_ | _0432_;
  assign _0434_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][7] [1] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][3] [1];
  assign _0633_ = ~ _0434_;
  assign _0435_ = _0210_ & _0633_;
  assign _0634_ = _0207_ | _0435_;
  assign _0436_ = ~ _0634_;
  assign _0635_ = _0007_ | _0016_;
  assign _0636_ = _0433_ & _0436_;
  assign _0437_ = ~ _0636_;
  assign _0438_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][11] [1] | _0208_;
  assign _0439_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][15] [1] | _0985_;
  assign _0440_ = _0210_ & _0439_;
  assign \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_credit_receiver/credit_incr [0] = ~ _0635_;
  assign _0637_ = _0438_ & _0440_;
  assign _0441_ = ~ _0637_;
  assign _0442_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][14] [1] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][10] [1];
  assign _0638_ = ~ _0442_;
  assign _0443_ = _0210_ | _0638_;
  assign _0639_ = _0441_ & _0443_;
  assign _0444_ = ~ _0639_;
  assign _0640_ = _0207_ & _0444_;
  assign _0445_ = ~ _0640_;
  assign _0641_ = _0437_ & _0445_;
  assign _0446_ = ~ _0641_;
  assign _0447_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][13] [1] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][9] [1];
  assign \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_visible [3] = _0007_ ? \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_saved [3] : _0018_;
  assign _0448_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][5] [1] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][1] [1];
  assign _0449_ = _0207_ ? _0447_ : _0448_;
  assign _0450_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][12] [1] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][8] [1];
  assign _0451_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][4] [1] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][0] [1];
  assign _0452_ = _0207_ ? _0450_ : _0451_;
  assign _0453_ = _0210_ ? _0449_ : _0452_;
  assign _0454_ = _0209_ ? _0446_ : _0453_;
  assign pop_data[1] = _0206_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][16] [1] : _0454_;
  assign _0455_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][6] [0] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][2] [0];
  assign _0456_ = _0210_ | _0455_;
  assign \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_visible [2] = _0007_ ? \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_saved [2] : _0020_;
  assign _0457_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][7] [0] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][3] [0];
  assign _0642_ = ~ _0457_;
  assign _0458_ = _0210_ & _0642_;
  assign _0643_ = _0207_ | _0458_;
  assign _0459_ = ~ _0643_;
  assign _0644_ = _0456_ & _0459_;
  assign _0460_ = ~ _0644_;
  assign _0461_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][11] [0] | _0208_;
  assign _0462_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][15] [0] | _0985_;
  assign _0463_ = _0210_ & _0462_;
  assign _0645_ = _0461_ & _0463_;
  assign _0464_ = ~ _0645_;
  assign \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_visible [1] = _0007_ ? \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_saved [1] : _0022_;
  assign _0465_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][14] [0] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][10] [0];
  assign _0646_ = ~ _0465_;
  assign _0466_ = _0210_ | _0646_;
  assign _0647_ = _0464_ & _0466_;
  assign _0467_ = ~ _0647_;
  assign _0648_ = _0207_ & _0467_;
  assign _0468_ = ~ _0648_;
  assign _0649_ = _0460_ & _0468_;
  assign _0469_ = ~ _0649_;
  assign _0470_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][13] [0] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][9] [0];
  assign _0471_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][5] [0] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][1] [0];
  assign _0472_ = _0207_ ? _0470_ : _0471_;
  assign \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_visible [0] = _0007_ ? \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_saved [0] : _0026_;
  assign _0473_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][12] [0] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][8] [0];
  assign _0474_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][4] [0] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][0] [0];
  assign _0475_ = _0207_ ? _0473_ : _0474_;
  assign _0476_ = _0210_ ? _0472_ : _0475_;
  assign _0477_ = _0209_ ? _0469_ : _0476_;
  assign pop_data[0] = _0206_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][16] [0] : _0477_;
  assign pop_items[1] = _0217_ ^ _0218_;
  assign _0478_ = _0210_ & \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_fifo_pop_ctrl_core/ram_rd_addr_update ;
  assign _0479_ = _0209_ & _0478_;
  assign _0480_ = _0208_ & _0479_;
  assign _0481_ = _0207_ & _0480_;
  assign _0482_ = _0206_ | _0481_;
  assign _0197_ = _0207_ ^ _0480_;
  assign _0198_ = _0208_ ^ _0479_;
  assign _0650_ = _0210_ ^ \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_fifo_pop_ctrl_core/ram_rd_addr_update ;
  assign _0483_ = ~ _0650_;
  assign _0199_ = _0209_ ^ _0478_;
  assign _0651_ = ~ _0199_;
  assign _0484_ = _0483_ & _0651_;
  assign _0652_ = ~ _0198_;
  assign _0485_ = _0484_ & _0652_;
  assign _0653_ = ~ _0197_;
  assign _0486_ = _0485_ & _0653_;
  assign _0196_ = _0482_ & _0486_;
  assign _0654_ = _0482_ | _0483_;
  assign _0200_ = ~ _0654_;
  always_ff @(posedge push_clk)
    _0008_ <= _0001_;
  always_ff @(posedge pop_clk)
    _0048_ <= \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_bit_toggle_reset_active_push/src_bit_internal ;
  assign _0655_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/push_beat  ? _0488_ : _0493_;
  assign _0656_ = _0006_ ? 1'h0 : _0655_;
  always_ff @(posedge push_clk)
    _0493_ <= _0656_;
  assign _0657_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/push_beat  ? _0489_ : _0494_;
  assign _0658_ = _0006_ ? 1'h0 : _0657_;
  always_ff @(posedge push_clk)
    _0494_ <= _0658_;
  assign _0659_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/push_beat  ? _0490_ : _0495_;
  assign _0660_ = _0006_ ? 1'h0 : _0659_;
  always_ff @(posedge push_clk)
    _0495_ <= _0660_;
  assign _0661_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/push_beat  ? _0491_ : _0496_;
  assign _0662_ = _0006_ ? 1'h0 : _0661_;
  always_ff @(posedge push_clk)
    _0496_ <= _0662_;
  assign _0663_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/push_beat  ? _0492_ : _0497_;
  assign _0664_ = _0006_ ? 1'h0 : _0663_;
  always_ff @(posedge push_clk)
    _0497_ <= _0664_;
  assign _0498_ = ~ \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/push_beat ;
  always_ff @(posedge pop_clk)
    _0054_ <= _0048_;
  assign _0487_ = ~ _0493_;
  assign _0526_ = ~ _0494_;
  assign _0499_ = _0496_ & _0497_;
  assign _0515_ = _0495_ & _0499_;
  assign _0665_ = ~ _0497_;
  assign _0500_ = _0496_ & _0665_;
  assign _0513_ = _0495_ & _0500_;
  assign _0666_ = ~ _0496_;
  assign _0501_ = _0497_ & _0666_;
  assign _0511_ = _0495_ & _0501_;
  assign _0667_ = _0496_ | _0497_;
  assign _0502_ = ~ _0667_;
  assign _0510_ = _0495_ & _0502_;
  assign _0525_ = _0494_ & _0515_;
  assign _0524_ = _0494_ & _0513_;
  assign _0523_ = _0494_ & _0511_;
  always_ff @(posedge pop_clk)
    _0049_ <= \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_gray_count_sync_push2pop/gen_cdc_sync[0].br_cdc_bit_toggle_inst/src_bit_internal ;
  assign _0522_ = _0494_ & _0510_;
  assign _0668_ = ~ _0495_;
  assign _0516_ = _0499_ & _0668_;
  assign _0521_ = _0494_ & _0516_;
  assign _0514_ = _0500_ & _0668_;
  assign _0520_ = _0494_ & _0514_;
  assign _0512_ = _0501_ & _0668_;
  assign _0519_ = _0494_ & _0512_;
  assign _0503_ = _0502_ & _0668_;
  assign _0517_ = _0494_ & _0503_;
  assign _0518_ = _0526_ & _0503_;
  assign _0561_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/push_beat  & _0493_;
  assign _0504_ = ~ _0561_;
  assign _0669_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/push_beat  & _0497_;
  assign _0505_ = ~ _0669_;
  always_ff @(posedge pop_clk)
    _0055_ <= _0049_;
  assign _0670_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/push_beat  & _0499_;
  assign _0506_ = ~ _0670_;
  assign _0507_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/push_beat  & _0515_;
  assign _0508_ = _0494_ & _0507_;
  assign _0488_ = _0487_ ? _0508_ : _0498_;
  assign _0671_ = _0526_ ^ _0507_;
  assign _0489_ = ~ _0671_;
  assign _0672_ = _0495_ ^ _0506_;
  assign _0490_ = ~ _0672_;
  assign _0673_ = _0496_ ^ _0505_;
  assign _0491_ = ~ _0673_;
  assign _0509_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/push_beat  ^ _0497_;
  assign _0492_ = _0504_ & _0509_;
  assign _0674_ = pop_rst ? 1'h0 : _0527_;
  always_ff @(posedge pop_clk)
    _0528_ <= _0674_;
  always_ff @(posedge pop_clk)
    _0050_ <= \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_gray_count_sync_push2pop/gen_cdc_sync[1].br_cdc_bit_toggle_inst/src_bit_internal ;
  assign _0675_ = pop_rst ? 1'h0 : _0528_;
  always_ff @(posedge pop_clk)
    \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_gray_count_sync_pop2push/gen_cdc_sync[1].br_cdc_bit_toggle_inst/src_bit_internal  <= _0675_;
  assign _0676_ = pop_rst ? 1'h0 : _0529_;
  always_ff @(posedge pop_clk)
    _0530_ <= _0676_;
  assign _0677_ = pop_rst ? 1'h0 : _0530_;
  always_ff @(posedge pop_clk)
    \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_gray_count_sync_pop2push/gen_cdc_sync[2].br_cdc_bit_toggle_inst/src_bit_internal  <= _0677_;
  assign _0678_ = pop_rst ? 1'h0 : _0531_;
  always_ff @(posedge pop_clk)
    _0532_ <= _0678_;
  assign _0679_ = pop_rst ? 1'h0 : _0532_;
  always_ff @(posedge pop_clk)
    \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_gray_count_sync_pop2push/gen_cdc_sync[3].br_cdc_bit_toggle_inst/src_bit_internal  <= _0679_;
  assign _0680_ = pop_rst ? 1'h0 : _0195_;
  always_ff @(posedge pop_clk)
    _0533_ <= _0680_;
  always_ff @(posedge pop_clk)
    _0056_ <= _0050_;
  assign _0681_ = pop_rst ? 1'h0 : _0533_;
  always_ff @(posedge pop_clk)
    \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_gray_count_sync_pop2push/gen_cdc_sync[4].br_cdc_bit_toggle_inst/src_bit_internal  <= _0681_;
  assign _0682_ = pop_rst ? 1'h0 : \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_cdc_fifo_pop_flag_mgr/push_count_adjusted [4];
  always_ff @(posedge pop_clk)
    \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_cdc_fifo_pop_flag_mgr/push_count_saved [4] <= _0682_;
  assign _0683_ = pop_rst ? 1'h0 : \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_cdc_fifo_pop_flag_mgr/push_count_adjusted [3];
  always_ff @(posedge pop_clk)
    \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_cdc_fifo_pop_flag_mgr/push_count_saved [3] <= _0683_;
  assign _0684_ = pop_rst ? 1'h0 : \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_cdc_fifo_pop_flag_mgr/push_count_adjusted [2];
  always_ff @(posedge pop_clk)
    \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_cdc_fifo_pop_flag_mgr/push_count_saved [2] <= _0684_;
  assign _0685_ = pop_rst ? 1'h0 : \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_cdc_fifo_pop_flag_mgr/push_count_adjusted [1];
  always_ff @(posedge pop_clk)
    \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_cdc_fifo_pop_flag_mgr/push_count_saved [1] <= _0685_;
  assign _0686_ = pop_rst ? 1'h0 : \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_cdc_fifo_pop_flag_mgr/push_count_adjusted [0];
  always_ff @(posedge pop_clk)
    \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_cdc_fifo_pop_flag_mgr/push_count_saved [0] <= _0686_;
  always_ff @(posedge pop_clk)
    _0051_ <= \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_gray_count_sync_push2pop/gen_cdc_sync[2].br_cdc_bit_toggle_inst/src_bit_internal ;
  assign _0687_ = pop_rst ? 1'h0 : _0534_;
  always_ff @(posedge pop_clk)
    _0535_ <= _0687_;
  assign _0688_ = pop_rst ? 1'h0 : _0535_;
  always_ff @(posedge pop_clk)
    \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_gray_count_sync_pop2push/gen_cdc_sync[0].br_cdc_bit_toggle_inst/src_bit_internal  <= _0688_;
  assign _0527_ = _0202_ ^ _0203_;
  assign _0529_ = _0201_ ^ _0202_;
  assign _0531_ = _0195_ ^ _0201_;
  assign _0534_ = _0203_ ^ _0194_;
  assign _0689_ = _0536_ ? push_data[7] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][3] [7];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][3] [7] <= _0689_;
  assign _0690_ = _0536_ ? push_data[6] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][3] [6];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][3] [6] <= _0690_;
  assign _0691_ = _0536_ ? push_data[5] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][3] [5];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][3] [5] <= _0691_;
  assign _0692_ = _0536_ ? push_data[4] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][3] [4];
  always_ff @(posedge pop_clk)
    _0057_ <= _0051_;
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][3] [4] <= _0692_;
  assign _0693_ = _0536_ ? push_data[3] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][3] [3];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][3] [3] <= _0693_;
  assign _0694_ = _0536_ ? push_data[2] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][3] [2];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][3] [2] <= _0694_;
  assign _0695_ = _0536_ ? push_data[1] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][3] [1];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][3] [1] <= _0695_;
  assign _0696_ = _0536_ ? push_data[0] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][3] [0];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][3] [0] <= _0696_;
  assign _0537_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/push_beat  & _0487_;
  assign _0538_ = _0516_ & _0526_;
  assign _0536_ = _0537_ & _0538_;
  assign _0697_ = _0539_ ? push_data[7] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][2] [7];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][2] [7] <= _0697_;
  assign _0698_ = _0539_ ? push_data[6] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][2] [6];
  always_ff @(posedge pop_clk)
    _0052_ <= \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_gray_count_sync_push2pop/gen_cdc_sync[3].br_cdc_bit_toggle_inst/src_bit_internal ;
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][2] [6] <= _0698_;
  assign _0699_ = _0539_ ? push_data[5] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][2] [5];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][2] [5] <= _0699_;
  assign _0700_ = _0539_ ? push_data[4] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][2] [4];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][2] [4] <= _0700_;
  assign _0701_ = _0539_ ? push_data[3] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][2] [3];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][2] [3] <= _0701_;
  assign _0702_ = _0539_ ? push_data[2] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][2] [2];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][2] [2] <= _0702_;
  assign _0703_ = _0539_ ? push_data[1] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][2] [1];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][2] [1] <= _0703_;
  assign _0704_ = _0539_ ? push_data[0] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][2] [0];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][2] [0] <= _0704_;
  assign _0541_ = _0514_ & _0526_;
  assign _0539_ = _0537_ & _0541_;
  always_ff @(posedge pop_clk)
    _0058_ <= _0052_;
  assign _0705_ = _0542_ ? push_data[7] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][1] [7];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][1] [7] <= _0705_;
  assign _0706_ = _0542_ ? push_data[6] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][1] [6];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][1] [6] <= _0706_;
  assign _0707_ = _0542_ ? push_data[5] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][1] [5];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][1] [5] <= _0707_;
  assign _0708_ = _0542_ ? push_data[4] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][1] [4];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][1] [4] <= _0708_;
  assign _0709_ = _0542_ ? push_data[3] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][1] [3];
  always_ff @(posedge push_clk)
    _0002_ <= \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_gray_count_sync_pop2push/gen_cdc_sync[1].br_cdc_bit_toggle_inst/src_bit_internal ;
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][1] [3] <= _0709_;
  assign _0710_ = _0542_ ? push_data[2] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][1] [2];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][1] [2] <= _0710_;
  assign _0711_ = _0542_ ? push_data[1] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][1] [1];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][1] [1] <= _0711_;
  always_ff @(posedge pop_clk)
    _0053_ <= \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_gray_count_sync_push2pop/gen_cdc_sync[4].br_cdc_bit_toggle_inst/src_bit_internal ;
  assign _0712_ = _0542_ ? push_data[0] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][1] [0];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][1] [0] <= _0712_;
  assign _0544_ = _0512_ & _0526_;
  assign _0542_ = _0537_ & _0544_;
  assign _0713_ = _0545_ ? push_data[7] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][0] [7];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][0] [7] <= _0713_;
  assign _0714_ = _0545_ ? push_data[6] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][0] [6];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][0] [6] <= _0714_;
  assign _0715_ = _0545_ ? push_data[5] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][0] [5];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][0] [5] <= _0715_;
  assign _0716_ = _0545_ ? push_data[4] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][0] [4];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][0] [4] <= _0716_;
  assign _0717_ = _0545_ ? push_data[3] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][0] [3];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][0] [3] <= _0717_;
  always_ff @(posedge pop_clk)
    _0059_ <= _0053_;
  assign _0718_ = _0545_ ? push_data[2] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][0] [2];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][0] [2] <= _0718_;
  assign _0719_ = _0545_ ? push_data[1] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][0] [1];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][0] [1] <= _0719_;
  assign _0720_ = _0545_ ? push_data[0] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][0] [0];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][0] [0] <= _0720_;
  assign _0546_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/push_beat  & _0518_;
  assign _0545_ = _0487_ & _0546_;
  assign _0721_ = _0547_ ? push_data[7] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][14] [7];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][14] [7] <= _0721_;
  assign _0722_ = _0547_ ? push_data[6] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][14] [6];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][14] [6] <= _0722_;
  assign _0723_ = _0547_ ? push_data[5] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][14] [5];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][14] [5] <= _0723_;
  assign _0724_ = _0547_ ? push_data[4] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][14] [4];
  always_ff @(posedge pop_clk)
    \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_cdc_fifo_pop_flag_mgr/br_delay_nr_reset_active_pop/out_stages[1]  <= pop_rst;
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][14] [4] <= _0724_;
  assign _0725_ = _0547_ ? push_data[3] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][14] [3];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][14] [3] <= _0725_;
  assign _0726_ = _0547_ ? push_data[2] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][14] [2];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][14] [2] <= _0726_;
  assign \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_cdc_fifo_pop_flag_mgr/push_count_adjusted [4] = _0054_ ? \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_cdc_fifo_pop_flag_mgr/push_count_saved [4] : _0059_;
  assign _0727_ = _0547_ ? push_data[1] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][14] [1];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][14] [1] <= _0727_;
  assign _0728_ = _0547_ ? push_data[0] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][14] [0];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][14] [0] <= _0728_;
  assign _0548_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/push_beat  & _0524_;
  assign _0547_ = _0487_ & _0548_;
  assign _0729_ = _0549_ ? push_data[7] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][13] [7];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][13] [7] <= _0729_;
  assign _0730_ = _0549_ ? push_data[6] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][13] [6];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][13] [6] <= _0730_;
  assign _0060_ = _0058_ ^ _0059_;
  assign _0731_ = _0549_ ? push_data[5] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][13] [5];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][13] [5] <= _0731_;
  assign _0732_ = _0549_ ? push_data[4] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][13] [4];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][13] [4] <= _0732_;
  assign _0733_ = _0549_ ? push_data[3] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][13] [3];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][13] [3] <= _0733_;
  assign _0734_ = _0549_ ? push_data[2] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][13] [2];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][13] [2] <= _0734_;
  assign _0735_ = _0549_ ? push_data[1] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][13] [1];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][13] [1] <= _0735_;
  assign \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_cdc_fifo_pop_flag_mgr/push_count_adjusted [3] = _0054_ ? \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_cdc_fifo_pop_flag_mgr/push_count_saved [3] : _0060_;
  assign _0736_ = _0549_ ? push_data[0] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][13] [0];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][13] [0] <= _0736_;
  assign _0550_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/push_beat  & _0523_;
  assign _0549_ = _0487_ & _0550_;
  assign _0737_ = _0551_ ? push_data[7] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][12] [7];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][12] [7] <= _0737_;
  assign _0738_ = _0551_ ? push_data[6] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][12] [6];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][12] [6] <= _0738_;
  assign _0739_ = _0551_ ? push_data[5] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][12] [5];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][12] [5] <= _0739_;
  assign _0061_ = _0057_ ^ _0060_;
  assign _0740_ = _0551_ ? push_data[4] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][12] [4];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][12] [4] <= _0740_;
  assign _0741_ = _0551_ ? push_data[3] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][12] [3];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][12] [3] <= _0741_;
  assign _0742_ = _0551_ ? push_data[2] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][12] [2];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][12] [2] <= _0742_;
  assign _0743_ = _0551_ ? push_data[1] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][12] [1];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][12] [1] <= _0743_;
  assign _0744_ = _0551_ ? push_data[0] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][12] [0];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][12] [0] <= _0744_;
  assign _0552_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/push_beat  & _0522_;
  assign \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_cdc_fifo_pop_flag_mgr/push_count_adjusted [2] = _0054_ ? \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_cdc_fifo_pop_flag_mgr/push_count_saved [2] : _0061_;
  assign _0551_ = _0487_ & _0552_;
  assign _0745_ = _0553_ ? push_data[7] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][11] [7];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][11] [7] <= _0745_;
  assign _0746_ = _0553_ ? push_data[6] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][11] [6];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][11] [6] <= _0746_;
  assign _0747_ = _0553_ ? push_data[5] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][11] [5];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][11] [5] <= _0747_;
  assign _0748_ = _0553_ ? push_data[4] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][11] [4];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][11] [4] <= _0748_;
  assign _0062_ = _0056_ ^ _0061_;
  assign _0749_ = _0553_ ? push_data[3] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][11] [3];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][11] [3] <= _0749_;
  assign _0750_ = _0553_ ? push_data[2] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][11] [2];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][11] [2] <= _0750_;
  assign _0751_ = _0553_ ? push_data[1] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][11] [1];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][11] [1] <= _0751_;
  assign _0752_ = _0553_ ? push_data[0] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][11] [0];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][11] [0] <= _0752_;
  assign _0576_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/push_beat  & _0521_;
  assign _0553_ = _0487_ & _0554_;
  assign \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_cdc_fifo_pop_flag_mgr/push_count_adjusted [1] = _0054_ ? \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_cdc_fifo_pop_flag_mgr/push_count_saved [1] : _0062_;
  assign _0753_ = _0555_ ? push_data[7] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][10] [7];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][10] [7] <= _0753_;
  assign _0754_ = _0555_ ? push_data[6] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][10] [6];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][10] [6] <= _0754_;
  assign _0755_ = _0555_ ? push_data[5] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][10] [5];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][10] [5] <= _0755_;
  assign _0756_ = _0555_ ? push_data[4] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][10] [4];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][10] [4] <= _0756_;
  assign _0757_ = _0555_ ? push_data[3] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][10] [3];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][10] [3] <= _0757_;
  assign _0063_ = _0055_ ^ _0062_;
  assign _0758_ = _0555_ ? push_data[2] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][10] [2];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][10] [2] <= _0758_;
  assign _0759_ = _0555_ ? push_data[1] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][10] [1];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][10] [1] <= _0759_;
  assign _0760_ = _0555_ ? push_data[0] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][10] [0];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][10] [0] <= _0760_;
  assign _0556_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/push_beat  & _0520_;
  assign _0555_ = _0487_ & _0556_;
  assign _0761_ = _0557_ ? push_data[7] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][9] [7];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][9] [7] <= _0761_;
  assign \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_cdc_fifo_pop_flag_mgr/push_count_adjusted [0] = _0054_ ? \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_cdc_fifo_pop_flag_mgr/push_count_saved [0] : _0063_;
  assign _0762_ = _0557_ ? push_data[6] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][9] [6];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][9] [6] <= _0762_;
  assign _0763_ = _0557_ ? push_data[5] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][9] [5];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][9] [5] <= _0763_;
  assign _0764_ = _0557_ ? push_data[4] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][9] [4];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][9] [4] <= _0764_;
  assign _0765_ = _0557_ ? push_data[3] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][9] [3];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][9] [3] <= _0765_;
  assign _0766_ = _0557_ ? push_data[2] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][9] [2];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][9] [2] <= _0766_;
  assign _0767_ = _0557_ ? push_data[1] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][9] [1];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][9] [1] <= _0767_;
  assign _0768_ = _0557_ ? push_data[0] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][9] [0];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][9] [0] <= _0768_;
  assign _0558_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/push_beat  & _0519_;
  assign _0557_ = _0487_ & _0558_;
  assign _0769_ = _0559_ ? push_data[7] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][8] [7];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][8] [7] <= _0769_;
  assign _0770_ = _0559_ ? push_data[6] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][8] [6];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][8] [6] <= _0770_;
  assign _0771_ = _0559_ ? push_data[5] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][8] [5];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][8] [5] <= _0771_;
  assign _0772_ = _0559_ ? push_data[4] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][8] [4];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][8] [4] <= _0772_;
  assign _0773_ = _0559_ ? push_data[3] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][8] [3];
  assign _0774_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/push_beat  ? _0064_ : _0069_;
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][8] [3] <= _0773_;
  assign _0775_ = _0559_ ? push_data[2] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][8] [2];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][8] [2] <= _0775_;
  assign _0776_ = _0559_ ? push_data[1] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][8] [1];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][8] [1] <= _0776_;
  always_ff @(posedge push_clk)
    _0009_ <= _0002_;
  assign _0777_ = _0006_ ? 1'h0 : _0774_;
  assign _0778_ = _0559_ ? push_data[0] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][8] [0];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][8] [0] <= _0778_;
  assign _0560_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/push_beat  & _0517_;
  assign _0559_ = _0487_ & _0560_;
  assign _0779_ = _0561_ ? push_data[7] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][16] [7];
  always_ff @(posedge push_clk)
    _0069_ <= _0777_;
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][16] [7] <= _0779_;
  assign _0780_ = _0561_ ? push_data[6] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][16] [6];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][16] [6] <= _0780_;
  assign _0781_ = _0561_ ? push_data[5] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][16] [5];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][16] [5] <= _0781_;
  assign _0782_ = _0561_ ? push_data[4] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][16] [4];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][16] [4] <= _0782_;
  assign _0783_ = _0561_ ? push_data[3] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][16] [3];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][16] [3] <= _0783_;
  assign _0784_ = _0561_ ? push_data[2] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][16] [2];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][16] [2] <= _0784_;
  assign _0785_ = _0561_ ? push_data[1] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][16] [1];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][16] [1] <= _0785_;
  assign _0786_ = _0561_ ? push_data[0] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][16] [0];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][16] [0] <= _0786_;
  assign _0787_ = _0562_ ? push_data[7] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][7] [7];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][7] [7] <= _0787_;
  assign _0788_ = _0562_ ? push_data[6] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][7] [6];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][7] [6] <= _0788_;
  assign _0789_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/push_beat  ? _0065_ : _0070_;
  assign _0790_ = _0562_ ? push_data[5] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][7] [5];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][7] [5] <= _0790_;
  assign _0791_ = _0562_ ? push_data[4] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][7] [4];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][7] [4] <= _0791_;
  assign _0792_ = _0562_ ? push_data[3] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][7] [3];
  assign _0793_ = _0006_ ? 1'h0 : _0789_;
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][7] [3] <= _0792_;
  assign _0794_ = _0562_ ? push_data[2] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][7] [2];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][7] [2] <= _0794_;
  assign _0795_ = _0562_ ? push_data[1] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][7] [1];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][7] [1] <= _0795_;
  always_ff @(posedge push_clk)
    _0070_ <= _0793_;
  assign _0796_ = _0562_ ? push_data[0] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][7] [0];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][7] [0] <= _0796_;
  assign _0564_ = _0515_ & _0526_;
  assign _0562_ = _0537_ & _0564_;
  assign _0797_ = _0565_ ? push_data[7] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][6] [7];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][6] [7] <= _0797_;
  assign _0798_ = _0565_ ? push_data[6] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][6] [6];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][6] [6] <= _0798_;
  assign _0799_ = _0565_ ? push_data[5] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][6] [5];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][6] [5] <= _0799_;
  assign _0800_ = _0565_ ? push_data[4] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][6] [4];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][6] [4] <= _0800_;
  assign _0801_ = _0565_ ? push_data[3] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][6] [3];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][6] [3] <= _0801_;
  assign _0802_ = _0565_ ? push_data[2] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][6] [2];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][6] [2] <= _0802_;
  assign _0803_ = _0565_ ? push_data[1] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][6] [1];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][6] [1] <= _0803_;
  assign _0804_ = _0565_ ? push_data[0] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][6] [0];
  assign _0805_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/push_beat  ? _0066_ : _0071_;
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][6] [0] <= _0804_;
  assign _0567_ = _0513_ & _0526_;
  assign _0565_ = _0537_ & _0567_;
  assign _0806_ = _0568_ ? push_data[0] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][15] [0];
  assign _0807_ = _0006_ ? 1'h0 : _0805_;
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][15] [0] <= _0806_;
  assign _0808_ = _0568_ ? push_data[7] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][15] [7];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][15] [7] <= _0808_;
  assign _0809_ = _0568_ ? push_data[6] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][15] [6];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][15] [6] <= _0809_;
  always_ff @(posedge push_clk)
    _0071_ <= _0807_;
  assign _0810_ = _0568_ ? push_data[5] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][15] [5];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][15] [5] <= _0810_;
  assign _0811_ = _0568_ ? push_data[4] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][15] [4];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][15] [4] <= _0811_;
  assign _0812_ = _0568_ ? push_data[3] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][15] [3];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][15] [3] <= _0812_;
  assign _0813_ = _0568_ ? push_data[2] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][15] [2];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][15] [2] <= _0813_;
  assign _0814_ = _0568_ ? push_data[1] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][15] [1];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][15] [1] <= _0814_;
  assign _0569_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/push_beat  & _0525_;
  assign _0568_ = _0487_ & _0569_;
  assign _0815_ = _0570_ ? push_data[7] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][5] [7];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][5] [7] <= _0815_;
  assign _0816_ = _0570_ ? push_data[6] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][5] [6];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][5] [6] <= _0816_;
  assign _0817_ = _0570_ ? push_data[5] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][5] [5];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][5] [5] <= _0817_;
  assign _0818_ = _0570_ ? push_data[4] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][5] [4];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][5] [4] <= _0818_;
  assign _0819_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/push_beat  ? _0067_ : _0072_;
  assign _0820_ = _0570_ ? push_data[3] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][5] [3];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][5] [3] <= _0820_;
  assign _0821_ = _0570_ ? push_data[2] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][5] [2];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][5] [2] <= _0821_;
  assign _0822_ = _0570_ ? push_data[1] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][5] [1];
  assign _0823_ = _0006_ ? 1'h0 : _0819_;
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][5] [1] <= _0822_;
  assign _0824_ = _0570_ ? push_data[0] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][5] [0];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][5] [0] <= _0824_;
  assign _0572_ = _0511_ & _0526_;
  assign _0570_ = _0537_ & _0572_;
  always_ff @(posedge push_clk)
    _0072_ <= _0823_;
  assign _0825_ = _0573_ ? push_data[2] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][4] [2];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][4] [2] <= _0825_;
  assign _0826_ = _0573_ ? push_data[1] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][4] [1];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][4] [1] <= _0826_;
  assign _0827_ = _0573_ ? push_data[0] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][4] [0];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][4] [0] <= _0827_;
  assign _0828_ = _0573_ ? push_data[7] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][4] [7];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][4] [7] <= _0828_;
  assign _0829_ = _0573_ ? push_data[6] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][4] [6];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][4] [6] <= _0829_;
  assign _0830_ = _0573_ ? push_data[5] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][4] [5];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][4] [5] <= _0830_;
  assign _0831_ = _0573_ ? push_data[4] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][4] [4];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][4] [4] <= _0831_;
  assign _0832_ = _0573_ ? push_data[3] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][4] [3];
  always_ff @(posedge push_clk)
    \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][4] [3] <= _0832_;
  assign _0575_ = _0510_ & _0526_;
  assign _0573_ = _0537_ & _0575_;
  assign _0833_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/push_beat  ? _0068_ : _0073_;
  assign _0834_ = _0006_ ? 1'h0 : _0833_;
  always_ff @(posedge push_clk)
    _0073_ <= _0834_;
  assign _0100_ = ~ _0006_;
  assign _0835_ = ~ \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_visible [0];
  assign _0074_ = _0073_ | _0835_;
  always_ff @(posedge push_clk)
    _0003_ <= \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_gray_count_sync_pop2push/gen_cdc_sync[2].br_cdc_bit_toggle_inst/src_bit_internal ;
  assign _0836_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_visible [0] ^ _0073_;
  assign push_slots[0] = ~ _0836_;
  assign _0837_ = ~ _0072_;
  assign _0075_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_visible [1] | _0837_;
  assign _0838_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_visible [1] ^ _0072_;
  assign _0076_ = ~ _0838_;
  assign _0839_ = _0074_ & _0076_;
  assign _0077_ = ~ _0839_;
  assign _0840_ = _0075_ & _0077_;
  assign _0078_ = ~ _0840_;
  assign _0841_ = ~ _0071_;
  assign _0079_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_visible [2] | _0841_;
  assign _0842_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_visible [2] ^ _0071_;
  assign _0080_ = ~ _0842_;
  assign _0843_ = _0078_ & _0080_;
  assign _0081_ = ~ _0843_;
  assign _0844_ = _0078_ ^ _0080_;
  assign _0082_ = ~ _0844_;
  assign push_slots[1] = _0074_ ^ _0076_;
  always_ff @(posedge push_clk)
    _0010_ <= _0003_;
  assign _0845_ = ~ push_slots[1];
  assign _0083_ = _0082_ & _0845_;
  assign _0846_ = _0079_ & _0081_;
  assign _0084_ = ~ _0846_;
  assign _0847_ = ~ _0070_;
  assign _0085_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_visible [3] | _0847_;
  assign _0848_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_visible [3] ^ _0070_;
  assign _0086_ = ~ _0848_;
  assign _0849_ = _0084_ & _0086_;
  assign _0087_ = ~ _0849_;
  assign _0850_ = _0084_ ^ _0086_;
  assign _0088_ = ~ _0850_;
  assign _0089_ = _0083_ & _0088_;
  assign _0090_ = _0085_ & _0087_;
  assign _0851_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_visible [4] ^ _0069_;
  assign _0091_ = ~ _0851_;
  assign _0852_ = _0090_ ^ _0091_;
  assign _0092_ = ~ _0852_;
  assign _0853_ = _0089_ & _0092_;
  assign _0093_ = ~ _0853_;
  always_ff @(posedge push_clk)
    _0004_ <= \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_gray_count_sync_pop2push/gen_cdc_sync[3].br_cdc_bit_toggle_inst/src_bit_internal ;
  assign _0094_ = push_slots[0] | _0093_;
  assign push_full = ~ _0094_;
  assign _0095_ = push_valid & _0100_;
  assign \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/push_beat  = _0094_ & _0095_;
  assign _0096_ = _0073_ & \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/push_beat ;
  assign _0097_ = _0072_ & _0096_;
  assign _0098_ = _0071_ & _0097_;
  assign _0854_ = _0070_ & _0098_;
  assign _0099_ = ~ _0854_;
  assign _0855_ = _0069_ ^ _0099_;
  assign _0064_ = ~ _0855_;
  assign _0065_ = _0070_ ^ _0098_;
  assign _0066_ = _0071_ ^ _0097_;
  assign _0067_ = _0072_ ^ _0096_;
  assign _0068_ = _0073_ ^ \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/push_beat ;
  always_ff @(posedge push_clk)
    _0011_ <= _0004_;
  assign _0856_ = _0082_ ^ push_slots[1];
  assign push_slots[2] = ~ _0856_;
  assign push_slots[3] = _0083_ ^ _0088_;
  assign push_slots[4] = _0089_ ^ _0092_;
  assign _0857_ = _0006_ ? 1'h0 : \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_visible [4];
  always_ff @(posedge push_clk)
    \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_saved [4] <= _0857_;
  assign _0858_ = _0006_ ? 1'h0 : \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_visible [3];
  always_ff @(posedge push_clk)
    \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_saved [3] <= _0858_;
  always_ff @(posedge push_clk)
    _0005_ <= \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_gray_count_sync_pop2push/gen_cdc_sync[4].br_cdc_bit_toggle_inst/src_bit_internal ;
  assign _0859_ = _0006_ ? 1'h0 : \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_visible [2];
  always_ff @(posedge push_clk)
    \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_saved [2] <= _0859_;
  assign _0860_ = _0006_ ? 1'h0 : \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_visible [1];
  always_ff @(posedge push_clk)
    \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_saved [1] <= _0860_;
  assign _0861_ = _0006_ ? 1'h0 : \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_visible [0];
  always_ff @(posedge push_clk)
    \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_saved [0] <= _0861_;
  assign _0862_ = _0006_ ? 1'h0 : _0101_;
  always_ff @(posedge push_clk)
    _0102_ <= _0862_;
  assign _0863_ = _0006_ ? 1'h0 : _0102_;
  always_ff @(posedge push_clk)
    \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_gray_count_sync_push2pop/gen_cdc_sync[0].br_cdc_bit_toggle_inst/src_bit_internal  <= _0863_;
  assign _0864_ = _0006_ ? 1'h0 : _0103_;
  always_ff @(posedge push_clk)
    _0104_ <= _0864_;
  always_ff @(posedge push_clk)
    _0012_ <= _0005_;
  assign _0865_ = _0006_ ? 1'h0 : _0104_;
  always_ff @(posedge push_clk)
    \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_gray_count_sync_push2pop/gen_cdc_sync[1].br_cdc_bit_toggle_inst/src_bit_internal  <= _0865_;
  assign _0866_ = _0006_ ? 1'h0 : _0105_;
  always_ff @(posedge push_clk)
    _0106_ <= _0866_;
  assign _0867_ = _0006_ ? 1'h0 : _0106_;
  always_ff @(posedge push_clk)
    \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_gray_count_sync_push2pop/gen_cdc_sync[2].br_cdc_bit_toggle_inst/src_bit_internal  <= _0867_;
  assign _0868_ = _0006_ ? 1'h0 : _0107_;
  always_ff @(posedge push_clk)
    _0108_ <= _0868_;
  assign _0869_ = _0006_ ? 1'h0 : _0108_;
  always_ff @(posedge push_clk)
    \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_gray_count_sync_push2pop/gen_cdc_sync[3].br_cdc_bit_toggle_inst/src_bit_internal  <= _0869_;
  assign _0870_ = _0006_ ? 1'h0 : _0064_;
  always_ff @(posedge push_clk)
    _0109_ <= _0870_;
  always_ff @(posedge push_clk)
    \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_bit_toggle_reset_active_push/src_bit_internal  <= _0006_;
  assign _0871_ = _0006_ ? 1'h0 : _0109_;
  always_ff @(posedge push_clk)
    \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_gray_count_sync_push2pop/gen_cdc_sync[4].br_cdc_bit_toggle_inst/src_bit_internal  <= _0871_;
  assign _0047_ = ~ \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_saved [4];
  assign _0046_ = ~ \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_saved [3];
  assign _0045_ = ~ \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_saved [2];
  assign _0044_ = ~ \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_saved [1];
  assign _0006_ = push_rst | push_sender_in_reset;
  assign _0043_ = ~ \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_saved [0];
  assign _0101_ = _0067_ ^ _0068_;
  assign _0103_ = _0066_ ^ _0067_;
  assign _0105_ = _0065_ ^ _0066_;
  assign _0107_ = _0064_ ^ _0065_;
  assign _0872_ = _0110_ ? _0111_ : credit_count_push[4];
  always_ff @(posedge push_clk)
    credit_count_push[4] <= _0872_;
  assign _0873_ = _0110_ ? _0112_ : credit_count_push[3];
  always_ff @(posedge push_clk)
    credit_count_push[3] <= _0873_;
  assign \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_visible [4] = _0007_ ? \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_cdc_fifo_push_flag_mgr/pop_count_saved [4] : _0012_;
  assign _0874_ = _0110_ ? _0113_ : credit_count_push[2];
  always_ff @(posedge push_clk)
    credit_count_push[2] <= _0874_;
  assign _0875_ = _0110_ ? _0114_ : credit_count_push[1];
  always_ff @(posedge push_clk)
    credit_count_push[1] <= _0875_;
  assign _0876_ = _0110_ ? _0115_ : credit_count_push[0];
  always_ff @(posedge push_clk)
    credit_count_push[0] <= _0876_;
  assign _0142_ = ~ push_credit_stall;
  assign _0877_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_credit_receiver/credit_incr [3] & credit_count_push[3];
  assign _0143_ = ~ _0877_;
  assign _0878_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_credit_receiver/credit_incr [2] & credit_count_push[2];
  assign _0144_ = ~ _0878_;
  assign _0018_ = _0011_ ^ _0012_;
  assign _0879_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_credit_receiver/credit_incr [1] & credit_count_push[1];
  assign _0145_ = ~ _0879_;
  assign _0146_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_credit_receiver/credit_incr [0] & credit_count_push[0];
  assign _0147_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_credit_receiver/credit_incr [1] ^ credit_count_push[1];
  assign _0880_ = _0146_ & _0147_;
  assign _0148_ = ~ _0880_;
  assign _0017_ = ~ _0018_;
  assign _0881_ = _0145_ & _0148_;
  assign _0149_ = ~ _0881_;
  assign _0150_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_credit_receiver/credit_incr [2] ^ credit_count_push[2];
  assign _0882_ = _0149_ & _0150_;
  assign _0151_ = ~ _0882_;
  assign _0883_ = _0144_ & _0151_;
  assign _0152_ = ~ _0883_;
  assign _0153_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_credit_receiver/credit_incr [3] ^ credit_count_push[3];
  assign _0884_ = _0152_ & _0153_;
  assign _0154_ = ~ _0884_;
  assign _0155_ = _0143_ & _0154_;
  assign _0885_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_credit_receiver/credit_incr [4] ^ credit_count_push[4];
  assign _0156_ = ~ _0885_;
  assign _0886_ = _0155_ ^ _0156_;
  assign _0157_ = ~ _0886_;
  assign _0158_ = credit_withhold_push[4] | _0157_;
  assign _0887_ = credit_withhold_push[4] & _0157_;
  assign _0159_ = ~ _0887_;
  assign _0888_ = _0152_ ^ _0153_;
  assign _0160_ = ~ _0888_;
  assign _0889_ = credit_withhold_push[3] & _0160_;
  assign _0161_ = ~ _0889_;
  assign _0162_ = credit_withhold_push[3] | _0160_;
  assign _0890_ = _0149_ ^ _0150_;
  assign _0163_ = ~ _0890_;
  assign _0891_ = _0046_ & _0018_;
  assign _0892_ = credit_withhold_push[2] & _0163_;
  assign _0164_ = ~ _0892_;
  assign _0165_ = credit_withhold_push[2] | _0163_;
  assign _0893_ = _0146_ ^ _0147_;
  assign _0166_ = ~ _0893_;
  assign _0894_ = credit_withhold_push[1] & _0166_;
  assign _0019_ = ~ _0891_;
  assign _0167_ = ~ _0894_;
  assign _0168_ = credit_withhold_push[1] | _0166_;
  assign _0895_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_credit_receiver/credit_incr [0] ^ credit_count_push[0];
  assign _0169_ = ~ _0895_;
  assign _0170_ = credit_withhold_push[0] | _0169_;
  assign _0896_ = _0168_ & _0170_;
  assign _0171_ = ~ _0896_;
  assign _0897_ = _0167_ & _0171_;
  assign _0172_ = ~ _0897_;
  assign _0898_ = _0165_ & _0172_;
  assign _0173_ = ~ _0898_;
  assign _0174_ = _0164_ & _0173_;
  assign _0899_ = _0010_ ^ _0017_;
  assign _0900_ = _0161_ & _0174_;
  assign _0175_ = ~ _0900_;
  assign _0901_ = _0162_ & _0175_;
  assign _0176_ = ~ _0901_;
  assign _0902_ = _0159_ & _0176_;
  assign _0177_ = ~ _0902_;
  assign _0903_ = _0158_ & _0177_;
  assign _0020_ = ~ _0899_;
  assign _0178_ = ~ _0903_;
  assign _0179_ = _0142_ & _0178_;
  assign _0904_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_credit_receiver/credit_incr [2] | \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_credit_receiver/credit_incr [1];
  assign _0180_ = ~ _0904_;
  assign _0905_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_credit_receiver/credit_incr [4] | \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_credit_receiver/credit_incr [0];
  assign _0181_ = ~ _0905_;
  assign _0906_ = ~ \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_push_1r1w_push_credit_inst/br_cdc_fifo_push_ctrl_credit/br_credit_receiver/credit_incr [3];
  assign _0182_ = _0181_ & _0906_;
  assign _0907_ = _0180_ & _0182_;
  assign _0183_ = ~ _0907_;
  assign _0184_ = _0179_ | _0183_;
  assign _0110_ = _0006_ | _0184_;
  assign _0908_ = _0045_ & _0020_;
  assign _0185_ = _0161_ & _0162_;
  assign _0186_ = _0164_ & _0165_;
  assign _0187_ = _0167_ & _0168_;
  assign _0909_ = credit_withhold_push[0] & _0169_;
  assign _0188_ = ~ _0909_;
  assign _0910_ = _0187_ & _0188_;
  assign _0021_ = ~ _0908_;
  assign _0189_ = ~ _0910_;
  assign _0911_ = _0168_ & _0189_;
  assign _0190_ = ~ _0911_;
  assign _0912_ = _0186_ & _0190_;
  assign _0191_ = ~ _0912_;
  assign _0913_ = _0165_ & _0191_;
  assign _0192_ = ~ _0913_;
  always_ff @(posedge push_clk)
    _0000_ <= \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_cdc_fifo_pop_flag_mgr/br_delay_nr_reset_active_pop/out_stages[1] ;
  assign _0914_ = _0185_ & _0192_;
  assign _0193_ = ~ _0914_;
  assign _0915_ = _0162_ & _0193_;
  assign _0116_ = ~ _0915_;
  assign _0916_ = ~ _0158_;
  assign credit_available_push[4] = _0116_ & _0916_;
  assign _0022_ = _0009_ ^ _0020_;
  assign _0117_ = _0185_ ^ _0192_;
  assign credit_available_push[3] = _0178_ & _0117_;
  assign _0118_ = _0186_ ^ _0190_;
  assign credit_available_push[2] = _0178_ & _0118_;
  assign _0119_ = _0187_ ^ _0188_;
  assign credit_available_push[1] = _0178_ & _0119_;
  assign _0917_ = _0170_ & _0188_;
  assign _0120_ = ~ _0917_;
  assign credit_available_push[0] = _0178_ & _0120_;
  assign push_credit = _0100_ & _0179_;
  assign _0918_ = _0006_ & credit_initial_push[4];
  assign _0919_ = _0044_ & _0022_;
  assign _0121_ = ~ _0918_;
  assign _0122_ = _0169_ & _0179_;
  assign _0123_ = _0166_ & _0122_;
  assign _0124_ = _0163_ & _0123_;
  assign _0920_ = _0160_ & _0124_;
  assign _0125_ = ~ _0920_;
  assign _0023_ = ~ _0919_;
  assign _0126_ = _0100_ & _0184_;
  assign _0921_ = ~ _0157_;
  assign _0127_ = _0126_ & _0921_;
  assign _0922_ = _0125_ & _0127_;
  assign _0128_ = ~ _0922_;
  assign _0923_ = _0121_ & _0128_;
  assign _0111_ = ~ _0923_;
  assign _0924_ = _0160_ ^ _0124_;
  assign _0129_ = ~ _0924_;
  assign _0925_ = _0126_ & _0129_;
  assign _0130_ = ~ _0925_;
  assign _0926_ = _0006_ & credit_initial_push[3];
  assign _0131_ = ~ _0926_;
  assign _0927_ = _0044_ ^ _0022_;
  assign _0928_ = _0130_ & _0131_;
  assign _0112_ = ~ _0928_;
  assign _0929_ = _0163_ ^ _0123_;
  assign _0132_ = ~ _0929_;
  assign _0930_ = _0126_ & _0132_;
  assign _0133_ = ~ _0930_;
  assign _0024_ = ~ _0927_;
  assign _0931_ = _0006_ & credit_initial_push[2];
  assign _0134_ = ~ _0931_;
  assign _0932_ = _0133_ & _0134_;
  assign _0113_ = ~ _0932_;
  assign _0933_ = _0166_ ^ _0122_;
  assign _0135_ = ~ _0933_;
  assign _0934_ = _0126_ & _0135_;
  assign _0136_ = ~ _0934_;
  assign _0935_ = _0006_ & credit_initial_push[1];
  assign _0137_ = ~ _0935_;
  assign _0936_ = _0136_ & _0137_;
  assign _0114_ = ~ _0936_;
  assign _0937_ = _0169_ ^ _0179_;
  assign _0138_ = ~ _0937_;
  assign _0938_ = _0008_ ^ _0022_;
  assign _0939_ = _0126_ & _0138_;
  assign _0139_ = ~ _0939_;
  assign _0940_ = _0006_ & credit_initial_push[0];
  assign _0140_ = ~ _0940_;
  assign _0941_ = _0139_ & _0140_;
  assign _0115_ = ~ _0941_;
  assign _0025_ = ~ _0938_;
  assign _0942_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_fifo_pop_ctrl_core/ram_rd_addr_update  ? _0194_ : _0204_;
  assign _0943_ = pop_rst ? 1'h0 : _0942_;
  always_ff @(posedge pop_clk)
    _0204_ <= _0943_;
  assign _0944_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_fifo_pop_ctrl_core/ram_rd_addr_update  ? _0195_ : _0205_;
  assign _0945_ = pop_rst ? 1'h0 : _0944_;
  always_ff @(posedge pop_clk)
    _0205_ <= _0945_;
  assign _0946_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_fifo_pop_ctrl_core/ram_rd_addr_update  ? _0196_ : _0206_;
  assign _0947_ = pop_rst ? 1'h0 : _0946_;
  always_ff @(posedge pop_clk)
    _0206_ <= _0947_;
  assign _0026_ = ~ _0025_;
  assign _0948_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_fifo_pop_ctrl_core/ram_rd_addr_update  ? _0197_ : _0207_;
  assign _0949_ = pop_rst ? 1'h0 : _0948_;
  always_ff @(posedge pop_clk)
    _0207_ <= _0949_;
  assign _0950_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_fifo_pop_ctrl_core/ram_rd_addr_update  ? _0198_ : _0208_;
  assign _0951_ = pop_rst ? 1'h0 : _0950_;
  always_ff @(posedge pop_clk)
    _0208_ <= _0951_;
  assign _0952_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_fifo_pop_ctrl_core/ram_rd_addr_update  ? _0199_ : _0209_;
  assign _0953_ = pop_rst ? 1'h0 : _0952_;
  always_ff @(posedge pop_clk)
    _0209_ <= _0953_;
  assign _0954_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_fifo_pop_ctrl_core/ram_rd_addr_update  ? _0200_ : _0210_;
  assign _0955_ = ~ _0043_;
  assign _0956_ = pop_rst ? 1'h0 : _0954_;
  always_ff @(posedge pop_clk)
    _0210_ <= _0956_;
  assign _0957_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_fifo_pop_ctrl_core/ram_rd_addr_update  ? _0201_ : _0211_;
  assign _0958_ = pop_rst ? 1'h0 : _0957_;
  always_ff @(posedge pop_clk)
    _0211_ <= _0958_;
  assign _0027_ = _0025_ & _0955_;
  assign _0959_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_fifo_pop_ctrl_core/ram_rd_addr_update  ? _0202_ : _0212_;
  assign _0960_ = pop_rst ? 1'h0 : _0959_;
  always_ff @(posedge pop_clk)
    _0212_ <= _0960_;
  assign _0961_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_fifo_pop_ctrl_core/ram_rd_addr_update  ? _0203_ : _0213_;
  assign _0962_ = pop_rst ? 1'h0 : _0961_;
  always_ff @(posedge pop_clk)
    _0213_ <= _0962_;
  assign _0963_ = ~ \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_cdc_fifo_pop_flag_mgr/push_count_adjusted [3];
  assign _0214_ = _0211_ | _0963_;
  assign _0964_ = ~ \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_cdc_fifo_pop_flag_mgr/push_count_adjusted [2];
  assign _0215_ = _0212_ | _0964_;
  assign _0965_ = ~ \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_cdc_fifo_pop_flag_mgr/push_count_adjusted [1];
  assign _0216_ = _0213_ | _0965_;
  assign _0966_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_cdc_fifo_pop_flag_mgr/push_count_adjusted [1] ^ _0213_;
  assign _0028_ = _0024_ | _0027_;
  assign _0217_ = ~ _0966_;
  assign _0967_ = ~ _0204_;
  assign _0218_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_cdc_fifo_pop_flag_mgr/push_count_adjusted [0] | _0967_;
  assign _0968_ = _0217_ & _0218_;
  assign _0219_ = ~ _0968_;
  assign _0969_ = _0216_ & _0219_;
  assign _0220_ = ~ _0969_;
  assign _0970_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_cdc_fifo_pop_flag_mgr/push_count_adjusted [2] ^ _0212_;
  assign _0221_ = ~ _0970_;
  assign _0971_ = _0220_ & _0221_;
  assign _0222_ = ~ _0971_;
  assign _0972_ = _0215_ & _0222_;
  assign _0223_ = ~ _0972_;
  assign _0029_ = _0023_ & _0028_;
  assign _0973_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_cdc_fifo_pop_flag_mgr/push_count_adjusted [3] ^ _0211_;
  assign _0224_ = ~ _0973_;
  assign _0974_ = _0223_ & _0224_;
  assign _0225_ = ~ _0974_;
  assign _0975_ = _0214_ & _0225_;
  assign _0226_ = ~ _0975_;
  assign _0976_ = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_cdc_fifo_pop_flag_mgr/push_count_adjusted [4] ^ _0205_;
  assign _0227_ = ~ _0976_;
  assign _0977_ = _0226_ ^ _0227_;
  assign _0228_ = ~ _0977_;
  assign pop_items[4] = ~ _0228_;
  assign pop_items[3] = _0223_ ^ _0224_;
  assign pop_items[2] = _0220_ ^ _0221_;
  assign _0978_ = _0045_ ^ _0020_;
  assign pop_items[0] = \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_cdc_fifo_pop_flag_mgr/push_count_adjusted [0] ^ _0204_;
  assign _0979_ = ~ pop_items[0];
  assign _0229_ = _0217_ & _0979_;
  assign _0980_ = ~ pop_items[2];
  assign _0230_ = _0229_ & _0980_;
  assign _0981_ = ~ pop_items[3];
  assign _0030_ = ~ _0978_;
  assign _0231_ = _0230_ & _0981_;
  assign _0982_ = _0228_ & _0231_;
  assign pop_valid = ~ _0982_;
  assign pop_empty = ~ pop_valid;
  assign \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_fifo_pop_ctrl_core/ram_rd_addr_update  = pop_ready & pop_valid;
  assign _0232_ = _0204_ & \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_fifo_pop_ctrl_core/ram_rd_addr_update ;
  assign _0194_ = _0204_ ^ \br_cdc_fifo_ctrl_1r1w_push_credit/br_cdc_fifo_ctrl_pop_1r1w_inst/br_cdc_fifo_pop_ctrl/br_fifo_pop_ctrl_core/ram_rd_addr_update ;
  assign _0233_ = _0213_ & _0232_;
  assign _0234_ = _0212_ & _0233_;
  assign _0983_ = _0211_ & _0234_;
  assign _0235_ = ~ _0983_;
  assign _0031_ = _0029_ | _0030_;
  assign _0984_ = _0205_ ^ _0235_;
  assign _0195_ = ~ _0984_;
  assign _0201_ = _0211_ ^ _0234_;
  assign _0202_ = _0212_ ^ _0233_;
  assign _0203_ = _0213_ ^ _0232_;
  assign _0985_ = ~ _0208_;
  assign _0236_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][13] [7] | _0985_;
  assign _0237_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][9] [7] | _0208_;
  assign _0238_ = _0210_ & _0237_;
  assign _0986_ = _0236_ & _0238_;
  assign _0239_ = ~ _0986_;
  assign _0240_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][12] [7] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][8] [7];
  assign _0987_ = _0021_ & _0031_;
  assign _0988_ = ~ _0210_;
  assign _0241_ = _0240_ & _0988_;
  assign _0989_ = _0209_ | _0241_;
  assign _0242_ = ~ _0989_;
  assign _0990_ = _0239_ & _0242_;
  assign _0243_ = ~ _0990_;
  assign _0032_ = ~ _0987_;
  assign _0244_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][14] [7] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][10] [7];
  assign _0991_ = ~ _0244_;
  assign _0245_ = _0210_ | _0991_;
  assign _0246_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][15] [7] | _0985_;
  assign _0247_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][11] [7] | _0208_;
  assign _0248_ = _0210_ & _0247_;
  assign _0992_ = _0246_ & _0248_;
  assign _0249_ = ~ _0992_;
  assign _0250_ = _0245_ & _0249_;
  assign _0993_ = _0209_ & _0250_;
  assign _0251_ = ~ _0993_;
  assign _0994_ = _0046_ ^ _0017_;
  assign _0252_ = _0207_ & _0243_;
  assign _0995_ = _0251_ & _0252_;
  assign _0253_ = ~ _0995_;
  assign _0254_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][2] [7] | _0208_;
  assign _0996_ = ~ \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][6] [7];
  assign _0255_ = _0208_ & _0996_;
  always_ff @(posedge push_clk)
    _0007_ <= _0000_;
  assign _0033_ = ~ _0994_;
  assign _0997_ = _0210_ | _0255_;
  assign _0256_ = ~ _0997_;
  assign _0998_ = _0254_ & _0256_;
  assign _0257_ = ~ _0998_;
  assign _0258_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][7] [7] | _0985_;
  assign _0259_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][3] [7] | _0208_;
  assign _0260_ = _0210_ & _0259_;
  assign _0999_ = _0258_ & _0260_;
  assign _0261_ = ~ _0999_;
  assign _0262_ = _0257_ & _0261_;
  assign _0263_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][4] [7] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][0] [7];
  assign _1000_ = _0032_ & _0033_;
  assign _1001_ = ~ _0263_;
  assign _0264_ = _0210_ | _1001_;
  assign _0265_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][5] [7] | _0985_;
  assign _0266_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][1] [7] | _0208_;
  assign _0267_ = _0210_ & _0266_;
  assign _0034_ = ~ _1000_;
  assign _1002_ = _0265_ & _0267_;
  assign _0268_ = ~ _1002_;
  assign _0269_ = _0264_ & _0268_;
  assign _0270_ = _0209_ ? _0262_ : _0269_;
  assign _0271_ = _0207_ | _0270_;
  assign _1003_ = _0253_ & _0271_;
  assign _0272_ = ~ _1003_;
  assign pop_data[7] = _0206_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][16] [7] : _0272_;
  assign _0273_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][13] [6] | _0985_;
  assign _0274_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][9] [6] | _0208_;
  assign _0275_ = _0210_ & _0274_;
  assign _0035_ = _0019_ & _0034_;
  assign _1004_ = _0273_ & _0275_;
  assign _0276_ = ~ _1004_;
  assign _0277_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][12] [6] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][8] [6];
  assign _0278_ = _0277_ & _0988_;
  assign _1005_ = _0209_ | _0278_;
  assign _0279_ = ~ _1005_;
  assign _1006_ = _0276_ & _0279_;
  assign _0280_ = ~ _1006_;
  assign _0281_ = _0208_ ? \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][14] [6] : \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][10] [6];
  assign _1007_ = ~ _0281_;
  assign _0282_ = _0210_ | _1007_;
  assign _1008_ = _0047_ ^ _0012_;
  assign _0283_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][15] [6] | _0985_;
  assign _0284_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][11] [6] | _0208_;
  assign _0285_ = _0210_ & _0284_;
  assign _1009_ = _0283_ & _0285_;
  assign _0286_ = ~ _1009_;
  assign _0036_ = ~ _1008_;
  assign _0287_ = _0282_ & _0286_;
  assign _1010_ = _0209_ & _0287_;
  assign _0288_ = ~ _1010_;
  assign _0289_ = _0207_ & _0280_;
  assign _1011_ = _0288_ & _0289_;
  assign _0290_ = ~ _1011_;
  assign _0291_ = \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][2] [6] | _0208_;
  assign _1012_ = ~ \br_ram_flops/gen_row[0].gen_col[0].br_ram_flops_tile/gen_multi_entry.gen_read_port[0].gen_structured_read.br_mux_bin_structured_gates_inst/in_stages[0][6] [6];
  assign _0292_ = _0208_ & _1012_;
  assign _1013_ = _0210_ | _0292_;
  assign _0293_ = ~ _1013_;
  assign _1014_ = _0291_ & _0293_;
  assign _0294_ = ~ _1014_;
  assign push_receiver_in_reset = push_rst;
endmodule

module shift_right(out_valid, in, shift, fill, out);
  wire _101_;
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _053_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  input [4:0] fill;
  wire [4:0] fill;
  input [49:0] in;
  wire [49:0] in;
  output [49:0] out;
  wire [49:0] out;
  output out_valid;
  wire out_valid;
  input [2:0] shift;
  wire [2:0] shift;
  assign _003_ = shift[0] ? in[33] : in[28];
  assign _039_ = shift[1] ? fill[0] : _038_;
  assign out[45] = shift[2] ? fill[0] : _039_;
  assign _040_ = shift[0] ? in[49] : in[44];
  assign _041_ = shift[1] ? fill[4] : _040_;
  assign out[44] = shift[2] ? fill[4] : _041_;
  assign _042_ = shift[0] ? in[48] : in[43];
  assign _043_ = shift[1] ? fill[3] : _042_;
  assign out[43] = shift[2] ? fill[3] : _043_;
  assign _044_ = shift[0] ? in[47] : in[42];
  assign _045_ = shift[1] ? fill[2] : _044_;
  assign _004_ = shift[0] ? in[43] : in[38];
  assign out[42] = shift[2] ? fill[2] : _045_;
  assign _046_ = shift[0] ? in[46] : in[41];
  assign _047_ = shift[1] ? fill[1] : _046_;
  assign out[41] = shift[2] ? fill[1] : _047_;
  assign _048_ = shift[0] ? in[45] : in[40];
  assign _049_ = shift[1] ? fill[0] : _048_;
  assign out[40] = shift[2] ? fill[0] : _049_;
  assign _050_ = shift[0] ? in[44] : in[39];
  assign _051_ = shift[1] ? _024_ : _050_;
  assign out[39] = shift[2] ? fill[4] : _051_;
  assign _005_ = shift[1] ? _004_ : _003_;
  assign _053_ = shift[0] ? in[18] : in[13];
  assign _055_ = shift[0] ? in[28] : in[23];
  assign _056_ = shift[0] ? in[38] : in[33];
  assign _057_ = shift[1] ? _056_ : _055_;
  assign out[3] = shift[2] ? _057_ : 1'h0;
  assign _058_ = shift[1] ? _032_ : _004_;
  assign out[38] = shift[2] ? fill[3] : _058_;
  assign _059_ = shift[1] ? _034_ : _010_;
  assign out[8] = shift[2] ? _005_ : _002_;
  assign out[37] = shift[2] ? fill[2] : _059_;
  assign _060_ = shift[1] ? _036_ : _016_;
  assign out[36] = shift[2] ? fill[1] : _060_;
  assign _061_ = shift[1] ? _038_ : _022_;
  assign out[35] = shift[2] ? fill[0] : _061_;
  assign _062_ = shift[1] ? _040_ : _030_;
  assign out[34] = shift[2] ? fill[4] : _062_;
  assign _063_ = shift[1] ? _042_ : _056_;
  assign out[33] = shift[2] ? fill[3] : _063_;
  assign _064_ = shift[0] ? in[37] : in[32];
  assign _006_ = shift[0] ? in[12] : in[7];
  assign _065_ = shift[1] ? _044_ : _064_;
  assign out[32] = shift[2] ? fill[2] : _065_;
  assign _066_ = shift[0] ? in[36] : in[31];
  assign _067_ = shift[1] ? _046_ : _066_;
  assign out[31] = shift[2] ? fill[1] : _067_;
  assign _068_ = shift[0] ? in[35] : in[30];
  assign _069_ = shift[1] ? _048_ : _068_;
  assign out[30] = shift[2] ? fill[0] : _069_;
  assign _070_ = shift[0] ? in[34] : in[29];
  assign _071_ = shift[1] ? _050_ : _070_;
  assign _007_ = shift[0] ? in[22] : in[17];
  assign out[29] = shift[2] ? _025_ : _071_;
  assign _072_ = shift[0] ? in[7] : in[2];
  assign _073_ = shift[0] ? in[17] : in[12];
  assign _074_ = shift[1] ? _073_ : _072_;
  assign _075_ = shift[0] ? in[27] : in[22];
  assign _076_ = shift[1] ? _064_ : _075_;
  assign out[2] = shift[2] ? _076_ : _074_;
  assign out[28] = shift[2] ? _033_ : _005_;
  assign out[27] = shift[2] ? _035_ : _011_;
  assign out[26] = shift[2] ? _037_ : _017_;
  assign _008_ = shift[1] ? _007_ : _006_;
  assign out[25] = shift[2] ? _039_ : _023_;
  assign out[24] = shift[2] ? _041_ : _031_;
  assign out[23] = shift[2] ? _043_ : _057_;
  assign out[22] = shift[2] ? _045_ : _076_;
  assign _077_ = shift[0] ? in[26] : in[21];
  assign _078_ = shift[1] ? _066_ : _077_;
  assign out[21] = shift[2] ? _047_ : _078_;
  assign _079_ = shift[0] ? in[25] : in[20];
  assign _080_ = shift[1] ? _068_ : _079_;
  assign out[20] = shift[2] ? _049_ : _080_;
  assign _009_ = shift[0] ? in[32] : in[27];
  assign _081_ = shift[0] ? in[24] : in[19];
  assign _082_ = shift[1] ? _070_ : _081_;
  assign out[19] = shift[2] ? _051_ : _082_;
  assign _083_ = shift[0] ? in[6] : in[1];
  assign _084_ = shift[0] ? in[16] : in[11];
  assign _085_ = shift[1] ? _084_ : _083_;
  assign out[1] = shift[2] ? _078_ : _085_;
  assign _086_ = shift[1] ? _003_ : _001_;
  assign out[18] = shift[2] ? _058_ : _086_;
  assign _087_ = shift[1] ? _009_ : _007_;
  assign _010_ = shift[0] ? in[42] : in[37];
  assign out[17] = shift[2] ? _059_ : _087_;
  assign _088_ = shift[1] ? _015_ : _013_;
  assign out[16] = shift[2] ? _060_ : _088_;
  assign _089_ = shift[1] ? _021_ : _019_;
  assign out[15] = shift[2] ? _061_ : _089_;
  assign _090_ = shift[1] ? _029_ : _027_;
  assign out[14] = shift[2] ? _062_ : _090_;
  assign _091_ = shift[1] ? _055_ : _053_;
  assign out[13] = shift[2] ? _063_ : _091_;
  assign _092_ = shift[1] ? _075_ : _073_;
  assign _011_ = shift[1] ? _010_ : _009_;
  assign out[12] = shift[2] ? _065_ : _092_;
  assign _093_ = shift[1] ? _077_ : _084_;
  assign out[11] = shift[2] ? _067_ : _093_;
  assign _094_ = shift[0] ? in[15] : in[10];
  assign _095_ = shift[1] ? _079_ : _094_;
  assign out[10] = shift[2] ? _069_ : _095_;
  assign _096_ = shift[0] ? in[14] : in[9];
  assign _097_ = shift[1] ? _081_ : _096_;
  assign out[9] = shift[2] ? _071_ : _097_;
  assign _098_ = shift[0] ? in[5] : in[0];
  assign out[7] = shift[2] ? _011_ : _008_;
  assign _099_ = shift[1] ? _094_ : _098_;
  assign out[0] = shift[2] ? _080_ : _099_;
  assign _100_ = shift[1] | shift[0];
  assign _101_ = shift[2] & _100_;
  assign out_valid = ~ _101_;
  assign _012_ = shift[0] ? in[11] : in[6];
  assign _013_ = shift[0] ? in[21] : in[16];
  assign _014_ = shift[1] ? _013_ : _012_;
  assign _015_ = shift[0] ? in[31] : in[26];
  assign _000_ = shift[0] ? in[13] : in[8];
  assign _016_ = shift[0] ? in[41] : in[36];
  assign _017_ = shift[1] ? _016_ : _015_;
  assign out[6] = shift[2] ? _017_ : _014_;
  assign _018_ = shift[0] ? in[10] : in[5];
  assign _019_ = shift[0] ? in[20] : in[15];
  assign _020_ = shift[1] ? _019_ : _018_;
  assign _021_ = shift[0] ? in[30] : in[25];
  assign _022_ = shift[0] ? in[40] : in[35];
  assign _023_ = shift[1] ? _022_ : _021_;
  assign out[5] = shift[2] ? _023_ : _020_;
  assign _001_ = shift[0] ? in[23] : in[18];
  assign _024_ = shift[0] ? fill[4] : in[49];
  assign _025_ = shift[1] ? fill[4] : _024_;
  assign out[49] = shift[2] ? fill[4] : _025_;
  assign _026_ = shift[0] ? in[9] : in[4];
  assign _027_ = shift[0] ? in[19] : in[14];
  assign _028_ = shift[1] ? _027_ : _026_;
  assign _029_ = shift[0] ? in[29] : in[24];
  assign _030_ = shift[0] ? in[39] : in[34];
  assign _031_ = shift[1] ? _030_ : _029_;
  assign out[4] = shift[2] ? _031_ : _028_;
  assign _002_ = shift[1] ? _001_ : _000_;
  assign _032_ = shift[0] ? fill[3] : in[48];
  assign _033_ = shift[1] ? fill[3] : _032_;
  assign out[48] = shift[2] ? fill[3] : _033_;
  assign _034_ = shift[0] ? fill[2] : in[47];
  assign _035_ = shift[1] ? fill[2] : _034_;
  assign out[47] = shift[2] ? fill[2] : _035_;
  assign _036_ = shift[0] ? fill[1] : in[46];
  assign _037_ = shift[1] ? fill[1] : _036_;
  assign out[46] = shift[2] ? fill[1] : _037_;
  assign _038_ = shift[0] ? fill[0] : in[45];
endmodule

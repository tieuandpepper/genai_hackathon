module enc_bin2onehot(clk, rst, in_valid, in, out);
  wire _09_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  wire _08_;
  input clk;
  wire clk;
  input [3:0] in;
  wire [3:0] in;
  input in_valid;
  wire in_valid;
  output [14:0] out;
  wire [14:0] out;
  input rst;
  wire rst;
  assign _02_ = _01_ & _12_;
  assign out[1] = _00_ & _02_;
  assign _09_ = ~ in[0];
  assign _03_ = in_valid & _09_;
  assign _04_ = _03_ & _12_;
  assign out[0] = _00_ & _04_;
  assign _05_ = in[2] & in[3];
  assign _06_ = in[1] & _03_;
  assign out[14] = _05_ & _06_;
  assign out[13] = _02_ & _05_;
  assign out[12] = _04_ & _05_;
  assign _10_ = ~ in[2];
  assign _07_ = in[3] & _10_;
  assign _08_ = in[1] & _01_;
  assign out[11] = _07_ & _08_;
  assign out[10] = _06_ & _07_;
  assign _11_ = in[2] | in[3];
  assign out[9] = _02_ & _07_;
  assign out[8] = _04_ & _07_;
  assign _00_ = ~ _11_;
  assign out[3] = _00_ & _08_;
  assign out[2] = _00_ & _06_;
  assign _01_ = in_valid & in[0];
  assign _12_ = ~ in[1];
  assign out[7:4] = { _08_, _06_, _02_, _04_ };
endmodule
